// system_bd.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module system_bd (
		output wire        axi_ltc235x_cnv_if_pwm_0,                //    axi_ltc235x_cnv_if.pwm_0
		input  wire        axi_ltc235x_device_if_busy,              // axi_ltc235x_device_if.busy
		output wire        axi_ltc235x_device_if_lvds_cmos_n,       //                      .lvds_cmos_n
		output wire        axi_ltc235x_device_if_cs_n,              //                      .cs_n
		output wire        axi_ltc235x_device_if_pd,                //                      .pd
		output wire        axi_ltc235x_device_if_scki,              //                      .scki
		input  wire        axi_ltc235x_device_if_scko,              //                      .scko
		output wire        axi_ltc235x_device_if_sdi,               //                      .sdi
		input  wire        axi_ltc235x_device_if_sdo_0,             //                      .sdo_0
		input  wire        axi_ltc235x_device_if_sdo_1,             //                      .sdo_1
		input  wire        axi_ltc235x_device_if_sdo_2,             //                      .sdo_2
		input  wire        axi_ltc235x_device_if_sdo_3,             //                      .sdo_3
		input  wire        axi_ltc235x_device_if_sdo_4,             //                      .sdo_4
		input  wire        axi_ltc235x_device_if_sdo_5,             //                      .sdo_5
		input  wire        axi_ltc235x_device_if_sdo_6,             //                      .sdo_6
		input  wire        axi_ltc235x_device_if_sdo_7,             //                      .sdo_7
		input  wire [31:0] pr_rom_data_nc_rom_data,                 //        pr_rom_data_nc.rom_data
		input  wire        sys_clk_clk,                             //               sys_clk.clk
		input  wire [31:0] sys_gpio_bd_in_port,                     //           sys_gpio_bd.in_port
		output wire [31:0] sys_gpio_bd_out_port,                    //                      .out_port
		input  wire [31:0] sys_gpio_in_export,                      //           sys_gpio_in.export
		output wire [31:0] sys_gpio_out_export,                     //          sys_gpio_out.export
		output wire        sys_hps_h2f_reset_reset_n,               //     sys_hps_h2f_reset.reset_n
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TX_CLK, //        sys_hps_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TXD0,   //                      .hps_io_emac1_inst_TXD0
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TXD1,   //                      .hps_io_emac1_inst_TXD1
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TXD2,   //                      .hps_io_emac1_inst_TXD2
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TXD3,   //                      .hps_io_emac1_inst_TXD3
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RXD0,   //                      .hps_io_emac1_inst_RXD0
		inout  wire        sys_hps_hps_io_hps_io_emac1_inst_MDIO,   //                      .hps_io_emac1_inst_MDIO
		output wire        sys_hps_hps_io_hps_io_emac1_inst_MDC,    //                      .hps_io_emac1_inst_MDC
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RX_CTL, //                      .hps_io_emac1_inst_RX_CTL
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TX_CTL, //                      .hps_io_emac1_inst_TX_CTL
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RX_CLK, //                      .hps_io_emac1_inst_RX_CLK
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RXD1,   //                      .hps_io_emac1_inst_RXD1
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RXD2,   //                      .hps_io_emac1_inst_RXD2
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RXD3,   //                      .hps_io_emac1_inst_RXD3
		inout  wire        sys_hps_hps_io_hps_io_qspi_inst_IO0,     //                      .hps_io_qspi_inst_IO0
		inout  wire        sys_hps_hps_io_hps_io_qspi_inst_IO1,     //                      .hps_io_qspi_inst_IO1
		inout  wire        sys_hps_hps_io_hps_io_qspi_inst_IO2,     //                      .hps_io_qspi_inst_IO2
		inout  wire        sys_hps_hps_io_hps_io_qspi_inst_IO3,     //                      .hps_io_qspi_inst_IO3
		output wire        sys_hps_hps_io_hps_io_qspi_inst_SS0,     //                      .hps_io_qspi_inst_SS0
		output wire        sys_hps_hps_io_hps_io_qspi_inst_CLK,     //                      .hps_io_qspi_inst_CLK
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_CMD,     //                      .hps_io_sdio_inst_CMD
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_D0,      //                      .hps_io_sdio_inst_D0
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_D1,      //                      .hps_io_sdio_inst_D1
		output wire        sys_hps_hps_io_hps_io_sdio_inst_CLK,     //                      .hps_io_sdio_inst_CLK
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_D2,      //                      .hps_io_sdio_inst_D2
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_D3,      //                      .hps_io_sdio_inst_D3
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D0,      //                      .hps_io_usb1_inst_D0
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D1,      //                      .hps_io_usb1_inst_D1
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D2,      //                      .hps_io_usb1_inst_D2
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D3,      //                      .hps_io_usb1_inst_D3
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D4,      //                      .hps_io_usb1_inst_D4
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D5,      //                      .hps_io_usb1_inst_D5
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D6,      //                      .hps_io_usb1_inst_D6
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D7,      //                      .hps_io_usb1_inst_D7
		input  wire        sys_hps_hps_io_hps_io_usb1_inst_CLK,     //                      .hps_io_usb1_inst_CLK
		output wire        sys_hps_hps_io_hps_io_usb1_inst_STP,     //                      .hps_io_usb1_inst_STP
		input  wire        sys_hps_hps_io_hps_io_usb1_inst_DIR,     //                      .hps_io_usb1_inst_DIR
		input  wire        sys_hps_hps_io_hps_io_usb1_inst_NXT,     //                      .hps_io_usb1_inst_NXT
		output wire        sys_hps_hps_io_hps_io_spim1_inst_CLK,    //                      .hps_io_spim1_inst_CLK
		output wire        sys_hps_hps_io_hps_io_spim1_inst_MOSI,   //                      .hps_io_spim1_inst_MOSI
		input  wire        sys_hps_hps_io_hps_io_spim1_inst_MISO,   //                      .hps_io_spim1_inst_MISO
		output wire        sys_hps_hps_io_hps_io_spim1_inst_SS0,    //                      .hps_io_spim1_inst_SS0
		input  wire        sys_hps_hps_io_hps_io_uart0_inst_RX,     //                      .hps_io_uart0_inst_RX
		output wire        sys_hps_hps_io_hps_io_uart0_inst_TX,     //                      .hps_io_uart0_inst_TX
		output wire        sys_hps_i2c0_out_data,                   //          sys_hps_i2c0.out_data
		input  wire        sys_hps_i2c0_sda,                        //                      .sda
		output wire        sys_hps_i2c0_clk_clk,                    //      sys_hps_i2c0_clk.clk
		input  wire        sys_hps_i2c0_scl_in_clk,                 //   sys_hps_i2c0_scl_in.clk
		output wire [14:0] sys_hps_memory_mem_a,                    //        sys_hps_memory.mem_a
		output wire [2:0]  sys_hps_memory_mem_ba,                   //                      .mem_ba
		output wire        sys_hps_memory_mem_ck,                   //                      .mem_ck
		output wire        sys_hps_memory_mem_ck_n,                 //                      .mem_ck_n
		output wire        sys_hps_memory_mem_cke,                  //                      .mem_cke
		output wire        sys_hps_memory_mem_cs_n,                 //                      .mem_cs_n
		output wire        sys_hps_memory_mem_ras_n,                //                      .mem_ras_n
		output wire        sys_hps_memory_mem_cas_n,                //                      .mem_cas_n
		output wire        sys_hps_memory_mem_we_n,                 //                      .mem_we_n
		output wire        sys_hps_memory_mem_reset_n,              //                      .mem_reset_n
		inout  wire [31:0] sys_hps_memory_mem_dq,                   //                      .mem_dq
		inout  wire [3:0]  sys_hps_memory_mem_dqs,                  //                      .mem_dqs
		inout  wire [3:0]  sys_hps_memory_mem_dqs_n,                //                      .mem_dqs_n
		output wire        sys_hps_memory_mem_odt,                  //                      .mem_odt
		output wire [3:0]  sys_hps_memory_mem_dm,                   //                      .mem_dm
		input  wire        sys_hps_memory_oct_rzqin,                //                      .oct_rzqin
		input  wire        sys_rst_reset_n,                         //               sys_rst.reset_n
		input  wire        sys_spi_MISO,                            //               sys_spi.MISO
		output wire        sys_spi_MOSI,                            //                      .MOSI
		output wire        sys_spi_SCLK,                            //                      .SCLK
		output wire        sys_spi_SS_n,                            //                      .SS_n
		output wire        vga_out_vga_if_vga_clk,                  //        vga_out_vga_if.vga_clk
		output wire        vga_out_vga_if_vga_hsync,                //                      .vga_hsync
		output wire        vga_out_vga_if_vga_vsync,                //                      .vga_vsync
		output wire [7:0]  vga_out_vga_if_vga_red,                  //                      .vga_red
		output wire [7:0]  vga_out_vga_if_vga_green,                //                      .vga_green
		output wire [7:0]  vga_out_vga_if_vga_blue                  //                      .vga_blue
	);

	wire          video_dmac_m_axis_tvalid;                                               // video_dmac:m_axis_valid -> vga_out:vdma_valid
	wire          video_dmac_m_axis_tready;                                               // vga_out:vdma_ready -> video_dmac:m_axis_ready
	wire          video_dmac_m_axis_tlast;                                                // video_dmac:m_axis_last -> vga_out:vdma_end_of_frame
	wire   [63:0] video_dmac_m_axis_tdata;                                                // video_dmac:m_axis_data -> vga_out:vdma_data
	wire          sys_hps_h2f_user0_clock_clk;                                            // sys_hps:h2f_user0_clk -> [mm_interconnect_2:sys_dma_clk_clk_clk, rst_controller_003:clk, sys_hps:f2h_sdram1_clk, sys_hps:f2h_sdram2_clk]
	wire          pixel_clk_pll_outclk0_clk;                                              // pixel_clk_pll:outclk_0 -> vga_out:reference_clk
	wire          pixel_clk_pll_outclk1_clk;                                              // pixel_clk_pll:outclk_1 -> [mm_interconnect_3:pixel_clk_pll_outclk1_clk, rst_controller_001:clk, rst_controller_004:clk, sys_hps:f2h_sdram0_clk, vga_out:vdma_clk, video_dmac:m_axis_aclk, video_dmac:m_src_axi_aclk]
	wire          axi_ltc235x_adc_ch_0_valid;                                             // axi_ltc235x:adc_valid_0 -> util_adc_pack:fifo_wr_en_0
	wire   [31:0] axi_ltc235x_adc_ch_0_data;                                              // axi_ltc235x:adc_data_0 -> util_adc_pack:fifo_wr_data_0
	wire          axi_ltc235x_adc_ch_0_enable;                                            // axi_ltc235x:adc_enable_0 -> util_adc_pack:enable_0
	wire          axi_ltc235x_adc_ch_1_valid;                                             // axi_ltc235x:adc_valid_1 -> util_adc_pack:fifo_wr_en_1
	wire   [31:0] axi_ltc235x_adc_ch_1_data;                                              // axi_ltc235x:adc_data_1 -> util_adc_pack:fifo_wr_data_1
	wire          axi_ltc235x_adc_ch_1_enable;                                            // axi_ltc235x:adc_enable_1 -> util_adc_pack:enable_1
	wire          axi_ltc235x_adc_ch_2_valid;                                             // axi_ltc235x:adc_valid_2 -> util_adc_pack:fifo_wr_en_2
	wire   [31:0] axi_ltc235x_adc_ch_2_data;                                              // axi_ltc235x:adc_data_2 -> util_adc_pack:fifo_wr_data_2
	wire          axi_ltc235x_adc_ch_2_enable;                                            // axi_ltc235x:adc_enable_2 -> util_adc_pack:enable_2
	wire          axi_ltc235x_adc_ch_3_valid;                                             // axi_ltc235x:adc_valid_3 -> util_adc_pack:fifo_wr_en_3
	wire   [31:0] axi_ltc235x_adc_ch_3_data;                                              // axi_ltc235x:adc_data_3 -> util_adc_pack:fifo_wr_data_3
	wire          axi_ltc235x_adc_ch_3_enable;                                            // axi_ltc235x:adc_enable_3 -> util_adc_pack:enable_3
	wire          axi_ltc235x_adc_ch_4_valid;                                             // axi_ltc235x:adc_valid_4 -> util_adc_pack:fifo_wr_en_4
	wire   [31:0] axi_ltc235x_adc_ch_4_data;                                              // axi_ltc235x:adc_data_4 -> util_adc_pack:fifo_wr_data_4
	wire          axi_ltc235x_adc_ch_4_enable;                                            // axi_ltc235x:adc_enable_4 -> util_adc_pack:enable_4
	wire          axi_ltc235x_adc_ch_5_valid;                                             // axi_ltc235x:adc_valid_5 -> util_adc_pack:fifo_wr_en_5
	wire   [31:0] axi_ltc235x_adc_ch_5_data;                                              // axi_ltc235x:adc_data_5 -> util_adc_pack:fifo_wr_data_5
	wire          axi_ltc235x_adc_ch_5_enable;                                            // axi_ltc235x:adc_enable_5 -> util_adc_pack:enable_5
	wire          axi_ltc235x_adc_ch_6_valid;                                             // axi_ltc235x:adc_valid_6 -> util_adc_pack:fifo_wr_en_6
	wire   [31:0] axi_ltc235x_adc_ch_6_data;                                              // axi_ltc235x:adc_data_6 -> util_adc_pack:fifo_wr_data_6
	wire          axi_ltc235x_adc_ch_6_enable;                                            // axi_ltc235x:adc_enable_6 -> util_adc_pack:enable_6
	wire          axi_ltc235x_adc_ch_7_valid;                                             // axi_ltc235x:adc_valid_7 -> util_adc_pack:fifo_wr_en_7
	wire   [31:0] axi_ltc235x_adc_ch_7_data;                                              // axi_ltc235x:adc_data_7 -> util_adc_pack:fifo_wr_data_7
	wire          axi_ltc235x_adc_ch_7_enable;                                            // axi_ltc235x:adc_enable_7 -> util_adc_pack:enable_7
	wire          util_adc_pack_if_fifo_wr_overflow_ovf;                                  // util_adc_pack:fifo_wr_overflow -> axi_ltc235x:adc_dovf
	wire          axi_adc_dma_if_fifo_wr_overflow_ovf;                                    // axi_adc_dma:fifo_wr_overflow -> util_adc_pack:packed_fifo_wr_overflow
	wire  [255:0] util_adc_pack_if_packed_fifo_wr_data_data;                              // util_adc_pack:packed_fifo_wr_data -> axi_adc_dma:fifo_wr_din
	wire          util_adc_pack_if_packed_fifo_wr_en_valid;                               // util_adc_pack:packed_fifo_wr_en -> axi_adc_dma:fifo_wr_en
	wire          util_adc_pack_if_packed_fifo_wr_sync_sync;                              // util_adc_pack:packed_fifo_wr_sync -> axi_adc_dma:fifo_wr_sync
	wire    [8:0] axi_sysid_0_if_rom_addr_rom_addr;                                       // axi_sysid_0:rom_addr -> rom_sys_0:rom_addr
	wire   [31:0] rom_sys_0_if_rom_data_rom_data;                                         // rom_sys_0:rom_data -> axi_sysid_0:sys_rom_data
	wire   [63:0] pixel_clk_pll_reconfig_from_pll_reconfig_from_pll;                      // pixel_clk_pll:reconfig_from_pll -> pixel_clk_pll_reconfig:reconfig_from_pll
	wire   [63:0] pixel_clk_pll_reconfig_reconfig_to_pll_reconfig_to_pll;                 // pixel_clk_pll_reconfig:reconfig_to_pll -> pixel_clk_pll:reconfig_to_pll
	wire    [1:0] sys_hps_h2f_axi_master_awburst;                                         // sys_hps:h2f_AWBURST -> mm_interconnect_0:sys_hps_h2f_axi_master_awburst
	wire    [3:0] sys_hps_h2f_axi_master_arlen;                                           // sys_hps:h2f_ARLEN -> mm_interconnect_0:sys_hps_h2f_axi_master_arlen
	wire    [7:0] sys_hps_h2f_axi_master_wstrb;                                           // sys_hps:h2f_WSTRB -> mm_interconnect_0:sys_hps_h2f_axi_master_wstrb
	wire          sys_hps_h2f_axi_master_wready;                                          // mm_interconnect_0:sys_hps_h2f_axi_master_wready -> sys_hps:h2f_WREADY
	wire   [11:0] sys_hps_h2f_axi_master_rid;                                             // mm_interconnect_0:sys_hps_h2f_axi_master_rid -> sys_hps:h2f_RID
	wire          sys_hps_h2f_axi_master_rready;                                          // sys_hps:h2f_RREADY -> mm_interconnect_0:sys_hps_h2f_axi_master_rready
	wire    [3:0] sys_hps_h2f_axi_master_awlen;                                           // sys_hps:h2f_AWLEN -> mm_interconnect_0:sys_hps_h2f_axi_master_awlen
	wire   [11:0] sys_hps_h2f_axi_master_wid;                                             // sys_hps:h2f_WID -> mm_interconnect_0:sys_hps_h2f_axi_master_wid
	wire    [3:0] sys_hps_h2f_axi_master_arcache;                                         // sys_hps:h2f_ARCACHE -> mm_interconnect_0:sys_hps_h2f_axi_master_arcache
	wire          sys_hps_h2f_axi_master_wvalid;                                          // sys_hps:h2f_WVALID -> mm_interconnect_0:sys_hps_h2f_axi_master_wvalid
	wire   [29:0] sys_hps_h2f_axi_master_araddr;                                          // sys_hps:h2f_ARADDR -> mm_interconnect_0:sys_hps_h2f_axi_master_araddr
	wire    [2:0] sys_hps_h2f_axi_master_arprot;                                          // sys_hps:h2f_ARPROT -> mm_interconnect_0:sys_hps_h2f_axi_master_arprot
	wire    [2:0] sys_hps_h2f_axi_master_awprot;                                          // sys_hps:h2f_AWPROT -> mm_interconnect_0:sys_hps_h2f_axi_master_awprot
	wire   [63:0] sys_hps_h2f_axi_master_wdata;                                           // sys_hps:h2f_WDATA -> mm_interconnect_0:sys_hps_h2f_axi_master_wdata
	wire          sys_hps_h2f_axi_master_arvalid;                                         // sys_hps:h2f_ARVALID -> mm_interconnect_0:sys_hps_h2f_axi_master_arvalid
	wire    [3:0] sys_hps_h2f_axi_master_awcache;                                         // sys_hps:h2f_AWCACHE -> mm_interconnect_0:sys_hps_h2f_axi_master_awcache
	wire   [11:0] sys_hps_h2f_axi_master_arid;                                            // sys_hps:h2f_ARID -> mm_interconnect_0:sys_hps_h2f_axi_master_arid
	wire    [1:0] sys_hps_h2f_axi_master_arlock;                                          // sys_hps:h2f_ARLOCK -> mm_interconnect_0:sys_hps_h2f_axi_master_arlock
	wire    [1:0] sys_hps_h2f_axi_master_awlock;                                          // sys_hps:h2f_AWLOCK -> mm_interconnect_0:sys_hps_h2f_axi_master_awlock
	wire   [29:0] sys_hps_h2f_axi_master_awaddr;                                          // sys_hps:h2f_AWADDR -> mm_interconnect_0:sys_hps_h2f_axi_master_awaddr
	wire    [1:0] sys_hps_h2f_axi_master_bresp;                                           // mm_interconnect_0:sys_hps_h2f_axi_master_bresp -> sys_hps:h2f_BRESP
	wire          sys_hps_h2f_axi_master_arready;                                         // mm_interconnect_0:sys_hps_h2f_axi_master_arready -> sys_hps:h2f_ARREADY
	wire   [63:0] sys_hps_h2f_axi_master_rdata;                                           // mm_interconnect_0:sys_hps_h2f_axi_master_rdata -> sys_hps:h2f_RDATA
	wire          sys_hps_h2f_axi_master_awready;                                         // mm_interconnect_0:sys_hps_h2f_axi_master_awready -> sys_hps:h2f_AWREADY
	wire    [1:0] sys_hps_h2f_axi_master_arburst;                                         // sys_hps:h2f_ARBURST -> mm_interconnect_0:sys_hps_h2f_axi_master_arburst
	wire    [2:0] sys_hps_h2f_axi_master_arsize;                                          // sys_hps:h2f_ARSIZE -> mm_interconnect_0:sys_hps_h2f_axi_master_arsize
	wire          sys_hps_h2f_axi_master_bready;                                          // sys_hps:h2f_BREADY -> mm_interconnect_0:sys_hps_h2f_axi_master_bready
	wire          sys_hps_h2f_axi_master_rlast;                                           // mm_interconnect_0:sys_hps_h2f_axi_master_rlast -> sys_hps:h2f_RLAST
	wire          sys_hps_h2f_axi_master_wlast;                                           // sys_hps:h2f_WLAST -> mm_interconnect_0:sys_hps_h2f_axi_master_wlast
	wire    [1:0] sys_hps_h2f_axi_master_rresp;                                           // mm_interconnect_0:sys_hps_h2f_axi_master_rresp -> sys_hps:h2f_RRESP
	wire   [11:0] sys_hps_h2f_axi_master_awid;                                            // sys_hps:h2f_AWID -> mm_interconnect_0:sys_hps_h2f_axi_master_awid
	wire   [11:0] sys_hps_h2f_axi_master_bid;                                             // mm_interconnect_0:sys_hps_h2f_axi_master_bid -> sys_hps:h2f_BID
	wire          sys_hps_h2f_axi_master_bvalid;                                          // mm_interconnect_0:sys_hps_h2f_axi_master_bvalid -> sys_hps:h2f_BVALID
	wire    [2:0] sys_hps_h2f_axi_master_awsize;                                          // sys_hps:h2f_AWSIZE -> mm_interconnect_0:sys_hps_h2f_axi_master_awsize
	wire          sys_hps_h2f_axi_master_awvalid;                                         // sys_hps:h2f_AWVALID -> mm_interconnect_0:sys_hps_h2f_axi_master_awvalid
	wire          sys_hps_h2f_axi_master_rvalid;                                          // mm_interconnect_0:sys_hps_h2f_axi_master_rvalid -> sys_hps:h2f_RVALID
	wire          mm_interconnect_0_sys_int_mem_s1_chipselect;                            // mm_interconnect_0:sys_int_mem_s1_chipselect -> sys_int_mem:chipselect
	wire   [63:0] mm_interconnect_0_sys_int_mem_s1_readdata;                              // sys_int_mem:readdata -> mm_interconnect_0:sys_int_mem_s1_readdata
	wire   [12:0] mm_interconnect_0_sys_int_mem_s1_address;                               // mm_interconnect_0:sys_int_mem_s1_address -> sys_int_mem:address
	wire    [7:0] mm_interconnect_0_sys_int_mem_s1_byteenable;                            // mm_interconnect_0:sys_int_mem_s1_byteenable -> sys_int_mem:byteenable
	wire          mm_interconnect_0_sys_int_mem_s1_write;                                 // mm_interconnect_0:sys_int_mem_s1_write -> sys_int_mem:write
	wire   [63:0] mm_interconnect_0_sys_int_mem_s1_writedata;                             // mm_interconnect_0:sys_int_mem_s1_writedata -> sys_int_mem:writedata
	wire          mm_interconnect_0_sys_int_mem_s1_clken;                                 // mm_interconnect_0:sys_int_mem_s1_clken -> sys_int_mem:clken
	wire    [1:0] sys_hps_h2f_lw_axi_master_awburst;                                      // sys_hps:h2f_lw_AWBURST -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_awburst
	wire    [3:0] sys_hps_h2f_lw_axi_master_arlen;                                        // sys_hps:h2f_lw_ARLEN -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_arlen
	wire    [3:0] sys_hps_h2f_lw_axi_master_wstrb;                                        // sys_hps:h2f_lw_WSTRB -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_wstrb
	wire          sys_hps_h2f_lw_axi_master_wready;                                       // mm_interconnect_1:sys_hps_h2f_lw_axi_master_wready -> sys_hps:h2f_lw_WREADY
	wire   [11:0] sys_hps_h2f_lw_axi_master_rid;                                          // mm_interconnect_1:sys_hps_h2f_lw_axi_master_rid -> sys_hps:h2f_lw_RID
	wire          sys_hps_h2f_lw_axi_master_rready;                                       // sys_hps:h2f_lw_RREADY -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_rready
	wire    [3:0] sys_hps_h2f_lw_axi_master_awlen;                                        // sys_hps:h2f_lw_AWLEN -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_awlen
	wire   [11:0] sys_hps_h2f_lw_axi_master_wid;                                          // sys_hps:h2f_lw_WID -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_wid
	wire    [3:0] sys_hps_h2f_lw_axi_master_arcache;                                      // sys_hps:h2f_lw_ARCACHE -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_arcache
	wire          sys_hps_h2f_lw_axi_master_wvalid;                                       // sys_hps:h2f_lw_WVALID -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_wvalid
	wire   [20:0] sys_hps_h2f_lw_axi_master_araddr;                                       // sys_hps:h2f_lw_ARADDR -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_araddr
	wire    [2:0] sys_hps_h2f_lw_axi_master_arprot;                                       // sys_hps:h2f_lw_ARPROT -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_arprot
	wire    [2:0] sys_hps_h2f_lw_axi_master_awprot;                                       // sys_hps:h2f_lw_AWPROT -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_awprot
	wire   [31:0] sys_hps_h2f_lw_axi_master_wdata;                                        // sys_hps:h2f_lw_WDATA -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_wdata
	wire          sys_hps_h2f_lw_axi_master_arvalid;                                      // sys_hps:h2f_lw_ARVALID -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_arvalid
	wire    [3:0] sys_hps_h2f_lw_axi_master_awcache;                                      // sys_hps:h2f_lw_AWCACHE -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_awcache
	wire   [11:0] sys_hps_h2f_lw_axi_master_arid;                                         // sys_hps:h2f_lw_ARID -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_arid
	wire    [1:0] sys_hps_h2f_lw_axi_master_arlock;                                       // sys_hps:h2f_lw_ARLOCK -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_arlock
	wire    [1:0] sys_hps_h2f_lw_axi_master_awlock;                                       // sys_hps:h2f_lw_AWLOCK -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_awlock
	wire   [20:0] sys_hps_h2f_lw_axi_master_awaddr;                                       // sys_hps:h2f_lw_AWADDR -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_awaddr
	wire    [1:0] sys_hps_h2f_lw_axi_master_bresp;                                        // mm_interconnect_1:sys_hps_h2f_lw_axi_master_bresp -> sys_hps:h2f_lw_BRESP
	wire          sys_hps_h2f_lw_axi_master_arready;                                      // mm_interconnect_1:sys_hps_h2f_lw_axi_master_arready -> sys_hps:h2f_lw_ARREADY
	wire   [31:0] sys_hps_h2f_lw_axi_master_rdata;                                        // mm_interconnect_1:sys_hps_h2f_lw_axi_master_rdata -> sys_hps:h2f_lw_RDATA
	wire          sys_hps_h2f_lw_axi_master_awready;                                      // mm_interconnect_1:sys_hps_h2f_lw_axi_master_awready -> sys_hps:h2f_lw_AWREADY
	wire    [1:0] sys_hps_h2f_lw_axi_master_arburst;                                      // sys_hps:h2f_lw_ARBURST -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_arburst
	wire    [2:0] sys_hps_h2f_lw_axi_master_arsize;                                       // sys_hps:h2f_lw_ARSIZE -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_arsize
	wire          sys_hps_h2f_lw_axi_master_bready;                                       // sys_hps:h2f_lw_BREADY -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_bready
	wire          sys_hps_h2f_lw_axi_master_rlast;                                        // mm_interconnect_1:sys_hps_h2f_lw_axi_master_rlast -> sys_hps:h2f_lw_RLAST
	wire          sys_hps_h2f_lw_axi_master_wlast;                                        // sys_hps:h2f_lw_WLAST -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_wlast
	wire    [1:0] sys_hps_h2f_lw_axi_master_rresp;                                        // mm_interconnect_1:sys_hps_h2f_lw_axi_master_rresp -> sys_hps:h2f_lw_RRESP
	wire   [11:0] sys_hps_h2f_lw_axi_master_awid;                                         // sys_hps:h2f_lw_AWID -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_awid
	wire   [11:0] sys_hps_h2f_lw_axi_master_bid;                                          // mm_interconnect_1:sys_hps_h2f_lw_axi_master_bid -> sys_hps:h2f_lw_BID
	wire          sys_hps_h2f_lw_axi_master_bvalid;                                       // mm_interconnect_1:sys_hps_h2f_lw_axi_master_bvalid -> sys_hps:h2f_lw_BVALID
	wire    [2:0] sys_hps_h2f_lw_axi_master_awsize;                                       // sys_hps:h2f_lw_AWSIZE -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_awsize
	wire          sys_hps_h2f_lw_axi_master_awvalid;                                      // sys_hps:h2f_lw_AWVALID -> mm_interconnect_1:sys_hps_h2f_lw_axi_master_awvalid
	wire          sys_hps_h2f_lw_axi_master_rvalid;                                       // mm_interconnect_1:sys_hps_h2f_lw_axi_master_rvalid -> sys_hps:h2f_lw_RVALID
	wire   [31:0] mm_interconnect_1_sys_id_control_slave_readdata;                        // sys_id:readdata -> mm_interconnect_1:sys_id_control_slave_readdata
	wire    [0:0] mm_interconnect_1_sys_id_control_slave_address;                         // mm_interconnect_1:sys_id_control_slave_address -> sys_id:address
	wire   [31:0] mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_readdata;    // pixel_clk_pll_reconfig:mgmt_readdata -> mm_interconnect_1:pixel_clk_pll_reconfig_mgmt_avalon_slave_readdata
	wire          mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_waitrequest; // pixel_clk_pll_reconfig:mgmt_waitrequest -> mm_interconnect_1:pixel_clk_pll_reconfig_mgmt_avalon_slave_waitrequest
	wire    [5:0] mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_address;     // mm_interconnect_1:pixel_clk_pll_reconfig_mgmt_avalon_slave_address -> pixel_clk_pll_reconfig:mgmt_address
	wire          mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_read;        // mm_interconnect_1:pixel_clk_pll_reconfig_mgmt_avalon_slave_read -> pixel_clk_pll_reconfig:mgmt_read
	wire          mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_write;       // mm_interconnect_1:pixel_clk_pll_reconfig_mgmt_avalon_slave_write -> pixel_clk_pll_reconfig:mgmt_write
	wire   [31:0] mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_writedata;   // mm_interconnect_1:pixel_clk_pll_reconfig_mgmt_avalon_slave_writedata -> pixel_clk_pll_reconfig:mgmt_writedata
	wire          mm_interconnect_1_sys_gpio_bd_s1_chipselect;                            // mm_interconnect_1:sys_gpio_bd_s1_chipselect -> sys_gpio_bd:chipselect
	wire   [31:0] mm_interconnect_1_sys_gpio_bd_s1_readdata;                              // sys_gpio_bd:readdata -> mm_interconnect_1:sys_gpio_bd_s1_readdata
	wire    [1:0] mm_interconnect_1_sys_gpio_bd_s1_address;                               // mm_interconnect_1:sys_gpio_bd_s1_address -> sys_gpio_bd:address
	wire          mm_interconnect_1_sys_gpio_bd_s1_write;                                 // mm_interconnect_1:sys_gpio_bd_s1_write -> sys_gpio_bd:write_n
	wire   [31:0] mm_interconnect_1_sys_gpio_bd_s1_writedata;                             // mm_interconnect_1:sys_gpio_bd_s1_writedata -> sys_gpio_bd:writedata
	wire          mm_interconnect_1_sys_gpio_in_s1_chipselect;                            // mm_interconnect_1:sys_gpio_in_s1_chipselect -> sys_gpio_in:chipselect
	wire   [31:0] mm_interconnect_1_sys_gpio_in_s1_readdata;                              // sys_gpio_in:readdata -> mm_interconnect_1:sys_gpio_in_s1_readdata
	wire    [1:0] mm_interconnect_1_sys_gpio_in_s1_address;                               // mm_interconnect_1:sys_gpio_in_s1_address -> sys_gpio_in:address
	wire          mm_interconnect_1_sys_gpio_in_s1_write;                                 // mm_interconnect_1:sys_gpio_in_s1_write -> sys_gpio_in:write_n
	wire   [31:0] mm_interconnect_1_sys_gpio_in_s1_writedata;                             // mm_interconnect_1:sys_gpio_in_s1_writedata -> sys_gpio_in:writedata
	wire          mm_interconnect_1_sys_gpio_out_s1_chipselect;                           // mm_interconnect_1:sys_gpio_out_s1_chipselect -> sys_gpio_out:chipselect
	wire   [31:0] mm_interconnect_1_sys_gpio_out_s1_readdata;                             // sys_gpio_out:readdata -> mm_interconnect_1:sys_gpio_out_s1_readdata
	wire    [1:0] mm_interconnect_1_sys_gpio_out_s1_address;                              // mm_interconnect_1:sys_gpio_out_s1_address -> sys_gpio_out:address
	wire          mm_interconnect_1_sys_gpio_out_s1_write;                                // mm_interconnect_1:sys_gpio_out_s1_write -> sys_gpio_out:write_n
	wire   [31:0] mm_interconnect_1_sys_gpio_out_s1_writedata;                            // mm_interconnect_1:sys_gpio_out_s1_writedata -> sys_gpio_out:writedata
	wire   [14:0] mm_interconnect_1_axi_sysid_0_s_axi_awaddr;                             // mm_interconnect_1:axi_sysid_0_s_axi_awaddr -> axi_sysid_0:s_axi_awaddr
	wire    [1:0] mm_interconnect_1_axi_sysid_0_s_axi_bresp;                              // axi_sysid_0:s_axi_bresp -> mm_interconnect_1:axi_sysid_0_s_axi_bresp
	wire          mm_interconnect_1_axi_sysid_0_s_axi_arready;                            // axi_sysid_0:s_axi_arready -> mm_interconnect_1:axi_sysid_0_s_axi_arready
	wire   [31:0] mm_interconnect_1_axi_sysid_0_s_axi_rdata;                              // axi_sysid_0:s_axi_rdata -> mm_interconnect_1:axi_sysid_0_s_axi_rdata
	wire    [3:0] mm_interconnect_1_axi_sysid_0_s_axi_wstrb;                              // mm_interconnect_1:axi_sysid_0_s_axi_wstrb -> axi_sysid_0:s_axi_wstrb
	wire          mm_interconnect_1_axi_sysid_0_s_axi_wready;                             // axi_sysid_0:s_axi_wready -> mm_interconnect_1:axi_sysid_0_s_axi_wready
	wire          mm_interconnect_1_axi_sysid_0_s_axi_awready;                            // axi_sysid_0:s_axi_awready -> mm_interconnect_1:axi_sysid_0_s_axi_awready
	wire          mm_interconnect_1_axi_sysid_0_s_axi_rready;                             // mm_interconnect_1:axi_sysid_0_s_axi_rready -> axi_sysid_0:s_axi_rready
	wire          mm_interconnect_1_axi_sysid_0_s_axi_bready;                             // mm_interconnect_1:axi_sysid_0_s_axi_bready -> axi_sysid_0:s_axi_bready
	wire          mm_interconnect_1_axi_sysid_0_s_axi_wvalid;                             // mm_interconnect_1:axi_sysid_0_s_axi_wvalid -> axi_sysid_0:s_axi_wvalid
	wire   [14:0] mm_interconnect_1_axi_sysid_0_s_axi_araddr;                             // mm_interconnect_1:axi_sysid_0_s_axi_araddr -> axi_sysid_0:s_axi_araddr
	wire    [2:0] mm_interconnect_1_axi_sysid_0_s_axi_arprot;                             // mm_interconnect_1:axi_sysid_0_s_axi_arprot -> axi_sysid_0:s_axi_arprot
	wire    [1:0] mm_interconnect_1_axi_sysid_0_s_axi_rresp;                              // axi_sysid_0:s_axi_rresp -> mm_interconnect_1:axi_sysid_0_s_axi_rresp
	wire    [2:0] mm_interconnect_1_axi_sysid_0_s_axi_awprot;                             // mm_interconnect_1:axi_sysid_0_s_axi_awprot -> axi_sysid_0:s_axi_awprot
	wire   [31:0] mm_interconnect_1_axi_sysid_0_s_axi_wdata;                              // mm_interconnect_1:axi_sysid_0_s_axi_wdata -> axi_sysid_0:s_axi_wdata
	wire          mm_interconnect_1_axi_sysid_0_s_axi_arvalid;                            // mm_interconnect_1:axi_sysid_0_s_axi_arvalid -> axi_sysid_0:s_axi_arvalid
	wire          mm_interconnect_1_axi_sysid_0_s_axi_bvalid;                             // axi_sysid_0:s_axi_bvalid -> mm_interconnect_1:axi_sysid_0_s_axi_bvalid
	wire          mm_interconnect_1_axi_sysid_0_s_axi_awvalid;                            // mm_interconnect_1:axi_sysid_0_s_axi_awvalid -> axi_sysid_0:s_axi_awvalid
	wire          mm_interconnect_1_axi_sysid_0_s_axi_rvalid;                             // axi_sysid_0:s_axi_rvalid -> mm_interconnect_1:axi_sysid_0_s_axi_rvalid
	wire   [10:0] mm_interconnect_1_video_dmac_s_axi_awaddr;                              // mm_interconnect_1:video_dmac_s_axi_awaddr -> video_dmac:s_axi_awaddr
	wire    [1:0] mm_interconnect_1_video_dmac_s_axi_bresp;                               // video_dmac:s_axi_bresp -> mm_interconnect_1:video_dmac_s_axi_bresp
	wire          mm_interconnect_1_video_dmac_s_axi_arready;                             // video_dmac:s_axi_arready -> mm_interconnect_1:video_dmac_s_axi_arready
	wire   [31:0] mm_interconnect_1_video_dmac_s_axi_rdata;                               // video_dmac:s_axi_rdata -> mm_interconnect_1:video_dmac_s_axi_rdata
	wire    [3:0] mm_interconnect_1_video_dmac_s_axi_wstrb;                               // mm_interconnect_1:video_dmac_s_axi_wstrb -> video_dmac:s_axi_wstrb
	wire          mm_interconnect_1_video_dmac_s_axi_wready;                              // video_dmac:s_axi_wready -> mm_interconnect_1:video_dmac_s_axi_wready
	wire          mm_interconnect_1_video_dmac_s_axi_awready;                             // video_dmac:s_axi_awready -> mm_interconnect_1:video_dmac_s_axi_awready
	wire          mm_interconnect_1_video_dmac_s_axi_rready;                              // mm_interconnect_1:video_dmac_s_axi_rready -> video_dmac:s_axi_rready
	wire          mm_interconnect_1_video_dmac_s_axi_bready;                              // mm_interconnect_1:video_dmac_s_axi_bready -> video_dmac:s_axi_bready
	wire          mm_interconnect_1_video_dmac_s_axi_wvalid;                              // mm_interconnect_1:video_dmac_s_axi_wvalid -> video_dmac:s_axi_wvalid
	wire   [10:0] mm_interconnect_1_video_dmac_s_axi_araddr;                              // mm_interconnect_1:video_dmac_s_axi_araddr -> video_dmac:s_axi_araddr
	wire    [2:0] mm_interconnect_1_video_dmac_s_axi_arprot;                              // mm_interconnect_1:video_dmac_s_axi_arprot -> video_dmac:s_axi_arprot
	wire    [1:0] mm_interconnect_1_video_dmac_s_axi_rresp;                               // video_dmac:s_axi_rresp -> mm_interconnect_1:video_dmac_s_axi_rresp
	wire    [2:0] mm_interconnect_1_video_dmac_s_axi_awprot;                              // mm_interconnect_1:video_dmac_s_axi_awprot -> video_dmac:s_axi_awprot
	wire   [31:0] mm_interconnect_1_video_dmac_s_axi_wdata;                               // mm_interconnect_1:video_dmac_s_axi_wdata -> video_dmac:s_axi_wdata
	wire          mm_interconnect_1_video_dmac_s_axi_arvalid;                             // mm_interconnect_1:video_dmac_s_axi_arvalid -> video_dmac:s_axi_arvalid
	wire          mm_interconnect_1_video_dmac_s_axi_bvalid;                              // video_dmac:s_axi_bvalid -> mm_interconnect_1:video_dmac_s_axi_bvalid
	wire          mm_interconnect_1_video_dmac_s_axi_awvalid;                             // mm_interconnect_1:video_dmac_s_axi_awvalid -> video_dmac:s_axi_awvalid
	wire          mm_interconnect_1_video_dmac_s_axi_rvalid;                              // video_dmac:s_axi_rvalid -> mm_interconnect_1:video_dmac_s_axi_rvalid
	wire   [15:0] mm_interconnect_1_vga_out_s_axi_awaddr;                                 // mm_interconnect_1:vga_out_s_axi_awaddr -> vga_out:s_axi_awaddr
	wire    [1:0] mm_interconnect_1_vga_out_s_axi_bresp;                                  // vga_out:s_axi_bresp -> mm_interconnect_1:vga_out_s_axi_bresp
	wire          mm_interconnect_1_vga_out_s_axi_arready;                                // vga_out:s_axi_arready -> mm_interconnect_1:vga_out_s_axi_arready
	wire   [31:0] mm_interconnect_1_vga_out_s_axi_rdata;                                  // vga_out:s_axi_rdata -> mm_interconnect_1:vga_out_s_axi_rdata
	wire    [3:0] mm_interconnect_1_vga_out_s_axi_wstrb;                                  // mm_interconnect_1:vga_out_s_axi_wstrb -> vga_out:s_axi_wstrb
	wire          mm_interconnect_1_vga_out_s_axi_wready;                                 // vga_out:s_axi_wready -> mm_interconnect_1:vga_out_s_axi_wready
	wire          mm_interconnect_1_vga_out_s_axi_awready;                                // vga_out:s_axi_awready -> mm_interconnect_1:vga_out_s_axi_awready
	wire          mm_interconnect_1_vga_out_s_axi_rready;                                 // mm_interconnect_1:vga_out_s_axi_rready -> vga_out:s_axi_rready
	wire          mm_interconnect_1_vga_out_s_axi_bready;                                 // mm_interconnect_1:vga_out_s_axi_bready -> vga_out:s_axi_bready
	wire          mm_interconnect_1_vga_out_s_axi_wvalid;                                 // mm_interconnect_1:vga_out_s_axi_wvalid -> vga_out:s_axi_wvalid
	wire   [15:0] mm_interconnect_1_vga_out_s_axi_araddr;                                 // mm_interconnect_1:vga_out_s_axi_araddr -> vga_out:s_axi_araddr
	wire    [2:0] mm_interconnect_1_vga_out_s_axi_arprot;                                 // mm_interconnect_1:vga_out_s_axi_arprot -> vga_out:s_axi_arprot
	wire    [1:0] mm_interconnect_1_vga_out_s_axi_rresp;                                  // vga_out:s_axi_rresp -> mm_interconnect_1:vga_out_s_axi_rresp
	wire    [2:0] mm_interconnect_1_vga_out_s_axi_awprot;                                 // mm_interconnect_1:vga_out_s_axi_awprot -> vga_out:s_axi_awprot
	wire   [31:0] mm_interconnect_1_vga_out_s_axi_wdata;                                  // mm_interconnect_1:vga_out_s_axi_wdata -> vga_out:s_axi_wdata
	wire          mm_interconnect_1_vga_out_s_axi_arvalid;                                // mm_interconnect_1:vga_out_s_axi_arvalid -> vga_out:s_axi_arvalid
	wire          mm_interconnect_1_vga_out_s_axi_bvalid;                                 // vga_out:s_axi_bvalid -> mm_interconnect_1:vga_out_s_axi_bvalid
	wire          mm_interconnect_1_vga_out_s_axi_awvalid;                                // mm_interconnect_1:vga_out_s_axi_awvalid -> vga_out:s_axi_awvalid
	wire          mm_interconnect_1_vga_out_s_axi_rvalid;                                 // vga_out:s_axi_rvalid -> mm_interconnect_1:vga_out_s_axi_rvalid
	wire   [15:0] mm_interconnect_1_axi_ltc235x_s_axi_awaddr;                             // mm_interconnect_1:axi_ltc235x_s_axi_awaddr -> axi_ltc235x:s_axi_awaddr
	wire    [1:0] mm_interconnect_1_axi_ltc235x_s_axi_bresp;                              // axi_ltc235x:s_axi_bresp -> mm_interconnect_1:axi_ltc235x_s_axi_bresp
	wire          mm_interconnect_1_axi_ltc235x_s_axi_arready;                            // axi_ltc235x:s_axi_arready -> mm_interconnect_1:axi_ltc235x_s_axi_arready
	wire   [31:0] mm_interconnect_1_axi_ltc235x_s_axi_rdata;                              // axi_ltc235x:s_axi_rdata -> mm_interconnect_1:axi_ltc235x_s_axi_rdata
	wire    [3:0] mm_interconnect_1_axi_ltc235x_s_axi_wstrb;                              // mm_interconnect_1:axi_ltc235x_s_axi_wstrb -> axi_ltc235x:s_axi_wstrb
	wire          mm_interconnect_1_axi_ltc235x_s_axi_wready;                             // axi_ltc235x:s_axi_wready -> mm_interconnect_1:axi_ltc235x_s_axi_wready
	wire          mm_interconnect_1_axi_ltc235x_s_axi_awready;                            // axi_ltc235x:s_axi_awready -> mm_interconnect_1:axi_ltc235x_s_axi_awready
	wire          mm_interconnect_1_axi_ltc235x_s_axi_rready;                             // mm_interconnect_1:axi_ltc235x_s_axi_rready -> axi_ltc235x:s_axi_rready
	wire          mm_interconnect_1_axi_ltc235x_s_axi_bready;                             // mm_interconnect_1:axi_ltc235x_s_axi_bready -> axi_ltc235x:s_axi_bready
	wire          mm_interconnect_1_axi_ltc235x_s_axi_wvalid;                             // mm_interconnect_1:axi_ltc235x_s_axi_wvalid -> axi_ltc235x:s_axi_wvalid
	wire   [15:0] mm_interconnect_1_axi_ltc235x_s_axi_araddr;                             // mm_interconnect_1:axi_ltc235x_s_axi_araddr -> axi_ltc235x:s_axi_araddr
	wire    [2:0] mm_interconnect_1_axi_ltc235x_s_axi_arprot;                             // mm_interconnect_1:axi_ltc235x_s_axi_arprot -> axi_ltc235x:s_axi_arprot
	wire    [1:0] mm_interconnect_1_axi_ltc235x_s_axi_rresp;                              // axi_ltc235x:s_axi_rresp -> mm_interconnect_1:axi_ltc235x_s_axi_rresp
	wire    [2:0] mm_interconnect_1_axi_ltc235x_s_axi_awprot;                             // mm_interconnect_1:axi_ltc235x_s_axi_awprot -> axi_ltc235x:s_axi_awprot
	wire   [31:0] mm_interconnect_1_axi_ltc235x_s_axi_wdata;                              // mm_interconnect_1:axi_ltc235x_s_axi_wdata -> axi_ltc235x:s_axi_wdata
	wire          mm_interconnect_1_axi_ltc235x_s_axi_arvalid;                            // mm_interconnect_1:axi_ltc235x_s_axi_arvalid -> axi_ltc235x:s_axi_arvalid
	wire          mm_interconnect_1_axi_ltc235x_s_axi_bvalid;                             // axi_ltc235x:s_axi_bvalid -> mm_interconnect_1:axi_ltc235x_s_axi_bvalid
	wire          mm_interconnect_1_axi_ltc235x_s_axi_awvalid;                            // mm_interconnect_1:axi_ltc235x_s_axi_awvalid -> axi_ltc235x:s_axi_awvalid
	wire          mm_interconnect_1_axi_ltc235x_s_axi_rvalid;                             // axi_ltc235x:s_axi_rvalid -> mm_interconnect_1:axi_ltc235x_s_axi_rvalid
	wire   [15:0] mm_interconnect_1_adc_pwm_gen_s_axi_awaddr;                             // mm_interconnect_1:adc_pwm_gen_s_axi_awaddr -> adc_pwm_gen:s_axi_awaddr
	wire    [1:0] mm_interconnect_1_adc_pwm_gen_s_axi_bresp;                              // adc_pwm_gen:s_axi_bresp -> mm_interconnect_1:adc_pwm_gen_s_axi_bresp
	wire          mm_interconnect_1_adc_pwm_gen_s_axi_arready;                            // adc_pwm_gen:s_axi_arready -> mm_interconnect_1:adc_pwm_gen_s_axi_arready
	wire   [31:0] mm_interconnect_1_adc_pwm_gen_s_axi_rdata;                              // adc_pwm_gen:s_axi_rdata -> mm_interconnect_1:adc_pwm_gen_s_axi_rdata
	wire    [3:0] mm_interconnect_1_adc_pwm_gen_s_axi_wstrb;                              // mm_interconnect_1:adc_pwm_gen_s_axi_wstrb -> adc_pwm_gen:s_axi_wstrb
	wire          mm_interconnect_1_adc_pwm_gen_s_axi_wready;                             // adc_pwm_gen:s_axi_wready -> mm_interconnect_1:adc_pwm_gen_s_axi_wready
	wire          mm_interconnect_1_adc_pwm_gen_s_axi_awready;                            // adc_pwm_gen:s_axi_awready -> mm_interconnect_1:adc_pwm_gen_s_axi_awready
	wire          mm_interconnect_1_adc_pwm_gen_s_axi_rready;                             // mm_interconnect_1:adc_pwm_gen_s_axi_rready -> adc_pwm_gen:s_axi_rready
	wire          mm_interconnect_1_adc_pwm_gen_s_axi_bready;                             // mm_interconnect_1:adc_pwm_gen_s_axi_bready -> adc_pwm_gen:s_axi_bready
	wire          mm_interconnect_1_adc_pwm_gen_s_axi_wvalid;                             // mm_interconnect_1:adc_pwm_gen_s_axi_wvalid -> adc_pwm_gen:s_axi_wvalid
	wire   [15:0] mm_interconnect_1_adc_pwm_gen_s_axi_araddr;                             // mm_interconnect_1:adc_pwm_gen_s_axi_araddr -> adc_pwm_gen:s_axi_araddr
	wire    [2:0] mm_interconnect_1_adc_pwm_gen_s_axi_arprot;                             // mm_interconnect_1:adc_pwm_gen_s_axi_arprot -> adc_pwm_gen:s_axi_arprot
	wire    [1:0] mm_interconnect_1_adc_pwm_gen_s_axi_rresp;                              // adc_pwm_gen:s_axi_rresp -> mm_interconnect_1:adc_pwm_gen_s_axi_rresp
	wire    [2:0] mm_interconnect_1_adc_pwm_gen_s_axi_awprot;                             // mm_interconnect_1:adc_pwm_gen_s_axi_awprot -> adc_pwm_gen:s_axi_awprot
	wire   [31:0] mm_interconnect_1_adc_pwm_gen_s_axi_wdata;                              // mm_interconnect_1:adc_pwm_gen_s_axi_wdata -> adc_pwm_gen:s_axi_wdata
	wire          mm_interconnect_1_adc_pwm_gen_s_axi_arvalid;                            // mm_interconnect_1:adc_pwm_gen_s_axi_arvalid -> adc_pwm_gen:s_axi_arvalid
	wire          mm_interconnect_1_adc_pwm_gen_s_axi_bvalid;                             // adc_pwm_gen:s_axi_bvalid -> mm_interconnect_1:adc_pwm_gen_s_axi_bvalid
	wire          mm_interconnect_1_adc_pwm_gen_s_axi_awvalid;                            // mm_interconnect_1:adc_pwm_gen_s_axi_awvalid -> adc_pwm_gen:s_axi_awvalid
	wire          mm_interconnect_1_adc_pwm_gen_s_axi_rvalid;                             // adc_pwm_gen:s_axi_rvalid -> mm_interconnect_1:adc_pwm_gen_s_axi_rvalid
	wire   [10:0] mm_interconnect_1_axi_adc_dma_s_axi_awaddr;                             // mm_interconnect_1:axi_adc_dma_s_axi_awaddr -> axi_adc_dma:s_axi_awaddr
	wire    [1:0] mm_interconnect_1_axi_adc_dma_s_axi_bresp;                              // axi_adc_dma:s_axi_bresp -> mm_interconnect_1:axi_adc_dma_s_axi_bresp
	wire          mm_interconnect_1_axi_adc_dma_s_axi_arready;                            // axi_adc_dma:s_axi_arready -> mm_interconnect_1:axi_adc_dma_s_axi_arready
	wire   [31:0] mm_interconnect_1_axi_adc_dma_s_axi_rdata;                              // axi_adc_dma:s_axi_rdata -> mm_interconnect_1:axi_adc_dma_s_axi_rdata
	wire    [3:0] mm_interconnect_1_axi_adc_dma_s_axi_wstrb;                              // mm_interconnect_1:axi_adc_dma_s_axi_wstrb -> axi_adc_dma:s_axi_wstrb
	wire          mm_interconnect_1_axi_adc_dma_s_axi_wready;                             // axi_adc_dma:s_axi_wready -> mm_interconnect_1:axi_adc_dma_s_axi_wready
	wire          mm_interconnect_1_axi_adc_dma_s_axi_awready;                            // axi_adc_dma:s_axi_awready -> mm_interconnect_1:axi_adc_dma_s_axi_awready
	wire          mm_interconnect_1_axi_adc_dma_s_axi_rready;                             // mm_interconnect_1:axi_adc_dma_s_axi_rready -> axi_adc_dma:s_axi_rready
	wire          mm_interconnect_1_axi_adc_dma_s_axi_bready;                             // mm_interconnect_1:axi_adc_dma_s_axi_bready -> axi_adc_dma:s_axi_bready
	wire          mm_interconnect_1_axi_adc_dma_s_axi_wvalid;                             // mm_interconnect_1:axi_adc_dma_s_axi_wvalid -> axi_adc_dma:s_axi_wvalid
	wire   [10:0] mm_interconnect_1_axi_adc_dma_s_axi_araddr;                             // mm_interconnect_1:axi_adc_dma_s_axi_araddr -> axi_adc_dma:s_axi_araddr
	wire    [2:0] mm_interconnect_1_axi_adc_dma_s_axi_arprot;                             // mm_interconnect_1:axi_adc_dma_s_axi_arprot -> axi_adc_dma:s_axi_arprot
	wire    [1:0] mm_interconnect_1_axi_adc_dma_s_axi_rresp;                              // axi_adc_dma:s_axi_rresp -> mm_interconnect_1:axi_adc_dma_s_axi_rresp
	wire    [2:0] mm_interconnect_1_axi_adc_dma_s_axi_awprot;                             // mm_interconnect_1:axi_adc_dma_s_axi_awprot -> axi_adc_dma:s_axi_awprot
	wire   [31:0] mm_interconnect_1_axi_adc_dma_s_axi_wdata;                              // mm_interconnect_1:axi_adc_dma_s_axi_wdata -> axi_adc_dma:s_axi_wdata
	wire          mm_interconnect_1_axi_adc_dma_s_axi_arvalid;                            // mm_interconnect_1:axi_adc_dma_s_axi_arvalid -> axi_adc_dma:s_axi_arvalid
	wire          mm_interconnect_1_axi_adc_dma_s_axi_bvalid;                             // axi_adc_dma:s_axi_bvalid -> mm_interconnect_1:axi_adc_dma_s_axi_bvalid
	wire          mm_interconnect_1_axi_adc_dma_s_axi_awvalid;                            // mm_interconnect_1:axi_adc_dma_s_axi_awvalid -> axi_adc_dma:s_axi_awvalid
	wire          mm_interconnect_1_axi_adc_dma_s_axi_rvalid;                             // axi_adc_dma:s_axi_rvalid -> mm_interconnect_1:axi_adc_dma_s_axi_rvalid
	wire          mm_interconnect_1_sys_spi_spi_control_port_chipselect;                  // mm_interconnect_1:sys_spi_spi_control_port_chipselect -> sys_spi:spi_select
	wire   [15:0] mm_interconnect_1_sys_spi_spi_control_port_readdata;                    // sys_spi:data_to_cpu -> mm_interconnect_1:sys_spi_spi_control_port_readdata
	wire    [2:0] mm_interconnect_1_sys_spi_spi_control_port_address;                     // mm_interconnect_1:sys_spi_spi_control_port_address -> sys_spi:mem_addr
	wire          mm_interconnect_1_sys_spi_spi_control_port_read;                        // mm_interconnect_1:sys_spi_spi_control_port_read -> sys_spi:read_n
	wire          mm_interconnect_1_sys_spi_spi_control_port_write;                       // mm_interconnect_1:sys_spi_spi_control_port_write -> sys_spi:write_n
	wire   [15:0] mm_interconnect_1_sys_spi_spi_control_port_writedata;                   // mm_interconnect_1:sys_spi_spi_control_port_writedata -> sys_spi:data_from_cpu
	wire    [1:0] axi_adc_dma_m_dest_axi_awburst;                                         // axi_adc_dma:m_dest_axi_awburst -> mm_interconnect_2:axi_adc_dma_m_dest_axi_awburst
	wire    [3:0] axi_adc_dma_m_dest_axi_arlen;                                           // axi_adc_dma:m_dest_axi_arlen -> mm_interconnect_2:axi_adc_dma_m_dest_axi_arlen
	wire    [7:0] axi_adc_dma_m_dest_axi_wstrb;                                           // axi_adc_dma:m_dest_axi_wstrb -> mm_interconnect_2:axi_adc_dma_m_dest_axi_wstrb
	wire          axi_adc_dma_m_dest_axi_wready;                                          // mm_interconnect_2:axi_adc_dma_m_dest_axi_wready -> axi_adc_dma:m_dest_axi_wready
	wire          axi_adc_dma_m_dest_axi_rid;                                             // mm_interconnect_2:axi_adc_dma_m_dest_axi_rid -> axi_adc_dma:m_dest_axi_rid
	wire          axi_adc_dma_m_dest_axi_rready;                                          // axi_adc_dma:m_dest_axi_rready -> mm_interconnect_2:axi_adc_dma_m_dest_axi_rready
	wire    [3:0] axi_adc_dma_m_dest_axi_awlen;                                           // axi_adc_dma:m_dest_axi_awlen -> mm_interconnect_2:axi_adc_dma_m_dest_axi_awlen
	wire          axi_adc_dma_m_dest_axi_wid;                                             // axi_adc_dma:m_dest_axi_wid -> mm_interconnect_2:axi_adc_dma_m_dest_axi_wid
	wire    [3:0] axi_adc_dma_m_dest_axi_arcache;                                         // axi_adc_dma:m_dest_axi_arcache -> mm_interconnect_2:axi_adc_dma_m_dest_axi_arcache
	wire          axi_adc_dma_m_dest_axi_wvalid;                                          // axi_adc_dma:m_dest_axi_wvalid -> mm_interconnect_2:axi_adc_dma_m_dest_axi_wvalid
	wire   [31:0] axi_adc_dma_m_dest_axi_araddr;                                          // axi_adc_dma:m_dest_axi_araddr -> mm_interconnect_2:axi_adc_dma_m_dest_axi_araddr
	wire    [2:0] axi_adc_dma_m_dest_axi_arprot;                                          // axi_adc_dma:m_dest_axi_arprot -> mm_interconnect_2:axi_adc_dma_m_dest_axi_arprot
	wire   [63:0] axi_adc_dma_m_dest_axi_wdata;                                           // axi_adc_dma:m_dest_axi_wdata -> mm_interconnect_2:axi_adc_dma_m_dest_axi_wdata
	wire          axi_adc_dma_m_dest_axi_arvalid;                                         // axi_adc_dma:m_dest_axi_arvalid -> mm_interconnect_2:axi_adc_dma_m_dest_axi_arvalid
	wire    [2:0] axi_adc_dma_m_dest_axi_awprot;                                          // axi_adc_dma:m_dest_axi_awprot -> mm_interconnect_2:axi_adc_dma_m_dest_axi_awprot
	wire    [3:0] axi_adc_dma_m_dest_axi_awcache;                                         // axi_adc_dma:m_dest_axi_awcache -> mm_interconnect_2:axi_adc_dma_m_dest_axi_awcache
	wire          axi_adc_dma_m_dest_axi_arid;                                            // axi_adc_dma:m_dest_axi_arid -> mm_interconnect_2:axi_adc_dma_m_dest_axi_arid
	wire    [1:0] axi_adc_dma_m_dest_axi_arlock;                                          // axi_adc_dma:m_dest_axi_arlock -> mm_interconnect_2:axi_adc_dma_m_dest_axi_arlock
	wire    [1:0] axi_adc_dma_m_dest_axi_awlock;                                          // axi_adc_dma:m_dest_axi_awlock -> mm_interconnect_2:axi_adc_dma_m_dest_axi_awlock
	wire   [31:0] axi_adc_dma_m_dest_axi_awaddr;                                          // axi_adc_dma:m_dest_axi_awaddr -> mm_interconnect_2:axi_adc_dma_m_dest_axi_awaddr
	wire    [1:0] axi_adc_dma_m_dest_axi_bresp;                                           // mm_interconnect_2:axi_adc_dma_m_dest_axi_bresp -> axi_adc_dma:m_dest_axi_bresp
	wire          axi_adc_dma_m_dest_axi_arready;                                         // mm_interconnect_2:axi_adc_dma_m_dest_axi_arready -> axi_adc_dma:m_dest_axi_arready
	wire   [63:0] axi_adc_dma_m_dest_axi_rdata;                                           // mm_interconnect_2:axi_adc_dma_m_dest_axi_rdata -> axi_adc_dma:m_dest_axi_rdata
	wire          axi_adc_dma_m_dest_axi_awready;                                         // mm_interconnect_2:axi_adc_dma_m_dest_axi_awready -> axi_adc_dma:m_dest_axi_awready
	wire    [1:0] axi_adc_dma_m_dest_axi_arburst;                                         // axi_adc_dma:m_dest_axi_arburst -> mm_interconnect_2:axi_adc_dma_m_dest_axi_arburst
	wire    [2:0] axi_adc_dma_m_dest_axi_arsize;                                          // axi_adc_dma:m_dest_axi_arsize -> mm_interconnect_2:axi_adc_dma_m_dest_axi_arsize
	wire          axi_adc_dma_m_dest_axi_bready;                                          // axi_adc_dma:m_dest_axi_bready -> mm_interconnect_2:axi_adc_dma_m_dest_axi_bready
	wire          axi_adc_dma_m_dest_axi_rlast;                                           // mm_interconnect_2:axi_adc_dma_m_dest_axi_rlast -> axi_adc_dma:m_dest_axi_rlast
	wire          axi_adc_dma_m_dest_axi_wlast;                                           // axi_adc_dma:m_dest_axi_wlast -> mm_interconnect_2:axi_adc_dma_m_dest_axi_wlast
	wire    [1:0] axi_adc_dma_m_dest_axi_rresp;                                           // mm_interconnect_2:axi_adc_dma_m_dest_axi_rresp -> axi_adc_dma:m_dest_axi_rresp
	wire          axi_adc_dma_m_dest_axi_awid;                                            // axi_adc_dma:m_dest_axi_awid -> mm_interconnect_2:axi_adc_dma_m_dest_axi_awid
	wire          axi_adc_dma_m_dest_axi_bid;                                             // mm_interconnect_2:axi_adc_dma_m_dest_axi_bid -> axi_adc_dma:m_dest_axi_bid
	wire          axi_adc_dma_m_dest_axi_bvalid;                                          // mm_interconnect_2:axi_adc_dma_m_dest_axi_bvalid -> axi_adc_dma:m_dest_axi_bvalid
	wire          axi_adc_dma_m_dest_axi_awvalid;                                         // axi_adc_dma:m_dest_axi_awvalid -> mm_interconnect_2:axi_adc_dma_m_dest_axi_awvalid
	wire          axi_adc_dma_m_dest_axi_rvalid;                                          // mm_interconnect_2:axi_adc_dma_m_dest_axi_rvalid -> axi_adc_dma:m_dest_axi_rvalid
	wire    [2:0] axi_adc_dma_m_dest_axi_awsize;                                          // axi_adc_dma:m_dest_axi_awsize -> mm_interconnect_2:axi_adc_dma_m_dest_axi_awsize
	wire    [1:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_awburst;                      // mm_interconnect_2:sys_hps_f2h_sdram1_data_awburst -> sys_hps:f2h_sdram1_AWBURST
	wire    [3:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_arlen;                        // mm_interconnect_2:sys_hps_f2h_sdram1_data_arlen -> sys_hps:f2h_sdram1_ARLEN
	wire    [7:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_wstrb;                        // mm_interconnect_2:sys_hps_f2h_sdram1_data_wstrb -> sys_hps:f2h_sdram1_WSTRB
	wire          mm_interconnect_2_sys_hps_f2h_sdram1_data_wready;                       // sys_hps:f2h_sdram1_WREADY -> mm_interconnect_2:sys_hps_f2h_sdram1_data_wready
	wire    [7:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_rid;                          // sys_hps:f2h_sdram1_RID -> mm_interconnect_2:sys_hps_f2h_sdram1_data_rid
	wire          mm_interconnect_2_sys_hps_f2h_sdram1_data_rready;                       // mm_interconnect_2:sys_hps_f2h_sdram1_data_rready -> sys_hps:f2h_sdram1_RREADY
	wire    [3:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_awlen;                        // mm_interconnect_2:sys_hps_f2h_sdram1_data_awlen -> sys_hps:f2h_sdram1_AWLEN
	wire    [7:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_wid;                          // mm_interconnect_2:sys_hps_f2h_sdram1_data_wid -> sys_hps:f2h_sdram1_WID
	wire    [3:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_arcache;                      // mm_interconnect_2:sys_hps_f2h_sdram1_data_arcache -> sys_hps:f2h_sdram1_ARCACHE
	wire          mm_interconnect_2_sys_hps_f2h_sdram1_data_wvalid;                       // mm_interconnect_2:sys_hps_f2h_sdram1_data_wvalid -> sys_hps:f2h_sdram1_WVALID
	wire   [31:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_araddr;                       // mm_interconnect_2:sys_hps_f2h_sdram1_data_araddr -> sys_hps:f2h_sdram1_ARADDR
	wire    [2:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_arprot;                       // mm_interconnect_2:sys_hps_f2h_sdram1_data_arprot -> sys_hps:f2h_sdram1_ARPROT
	wire    [2:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_awprot;                       // mm_interconnect_2:sys_hps_f2h_sdram1_data_awprot -> sys_hps:f2h_sdram1_AWPROT
	wire   [63:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_wdata;                        // mm_interconnect_2:sys_hps_f2h_sdram1_data_wdata -> sys_hps:f2h_sdram1_WDATA
	wire          mm_interconnect_2_sys_hps_f2h_sdram1_data_arvalid;                      // mm_interconnect_2:sys_hps_f2h_sdram1_data_arvalid -> sys_hps:f2h_sdram1_ARVALID
	wire    [3:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_awcache;                      // mm_interconnect_2:sys_hps_f2h_sdram1_data_awcache -> sys_hps:f2h_sdram1_AWCACHE
	wire    [7:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_arid;                         // mm_interconnect_2:sys_hps_f2h_sdram1_data_arid -> sys_hps:f2h_sdram1_ARID
	wire    [1:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_arlock;                       // mm_interconnect_2:sys_hps_f2h_sdram1_data_arlock -> sys_hps:f2h_sdram1_ARLOCK
	wire    [1:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_awlock;                       // mm_interconnect_2:sys_hps_f2h_sdram1_data_awlock -> sys_hps:f2h_sdram1_AWLOCK
	wire   [31:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_awaddr;                       // mm_interconnect_2:sys_hps_f2h_sdram1_data_awaddr -> sys_hps:f2h_sdram1_AWADDR
	wire    [1:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_bresp;                        // sys_hps:f2h_sdram1_BRESP -> mm_interconnect_2:sys_hps_f2h_sdram1_data_bresp
	wire          mm_interconnect_2_sys_hps_f2h_sdram1_data_arready;                      // sys_hps:f2h_sdram1_ARREADY -> mm_interconnect_2:sys_hps_f2h_sdram1_data_arready
	wire   [63:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_rdata;                        // sys_hps:f2h_sdram1_RDATA -> mm_interconnect_2:sys_hps_f2h_sdram1_data_rdata
	wire          mm_interconnect_2_sys_hps_f2h_sdram1_data_awready;                      // sys_hps:f2h_sdram1_AWREADY -> mm_interconnect_2:sys_hps_f2h_sdram1_data_awready
	wire    [1:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_arburst;                      // mm_interconnect_2:sys_hps_f2h_sdram1_data_arburst -> sys_hps:f2h_sdram1_ARBURST
	wire    [2:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_arsize;                       // mm_interconnect_2:sys_hps_f2h_sdram1_data_arsize -> sys_hps:f2h_sdram1_ARSIZE
	wire          mm_interconnect_2_sys_hps_f2h_sdram1_data_bready;                       // mm_interconnect_2:sys_hps_f2h_sdram1_data_bready -> sys_hps:f2h_sdram1_BREADY
	wire          mm_interconnect_2_sys_hps_f2h_sdram1_data_rlast;                        // sys_hps:f2h_sdram1_RLAST -> mm_interconnect_2:sys_hps_f2h_sdram1_data_rlast
	wire          mm_interconnect_2_sys_hps_f2h_sdram1_data_wlast;                        // mm_interconnect_2:sys_hps_f2h_sdram1_data_wlast -> sys_hps:f2h_sdram1_WLAST
	wire    [1:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_rresp;                        // sys_hps:f2h_sdram1_RRESP -> mm_interconnect_2:sys_hps_f2h_sdram1_data_rresp
	wire    [7:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_awid;                         // mm_interconnect_2:sys_hps_f2h_sdram1_data_awid -> sys_hps:f2h_sdram1_AWID
	wire    [7:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_bid;                          // sys_hps:f2h_sdram1_BID -> mm_interconnect_2:sys_hps_f2h_sdram1_data_bid
	wire          mm_interconnect_2_sys_hps_f2h_sdram1_data_bvalid;                       // sys_hps:f2h_sdram1_BVALID -> mm_interconnect_2:sys_hps_f2h_sdram1_data_bvalid
	wire    [2:0] mm_interconnect_2_sys_hps_f2h_sdram1_data_awsize;                       // mm_interconnect_2:sys_hps_f2h_sdram1_data_awsize -> sys_hps:f2h_sdram1_AWSIZE
	wire          mm_interconnect_2_sys_hps_f2h_sdram1_data_awvalid;                      // mm_interconnect_2:sys_hps_f2h_sdram1_data_awvalid -> sys_hps:f2h_sdram1_AWVALID
	wire          mm_interconnect_2_sys_hps_f2h_sdram1_data_rvalid;                       // sys_hps:f2h_sdram1_RVALID -> mm_interconnect_2:sys_hps_f2h_sdram1_data_rvalid
	wire    [1:0] video_dmac_m_src_axi_awburst;                                           // video_dmac:m_src_axi_awburst -> mm_interconnect_3:video_dmac_m_src_axi_awburst
	wire    [3:0] video_dmac_m_src_axi_arlen;                                             // video_dmac:m_src_axi_arlen -> mm_interconnect_3:video_dmac_m_src_axi_arlen
	wire    [7:0] video_dmac_m_src_axi_wstrb;                                             // video_dmac:m_src_axi_wstrb -> mm_interconnect_3:video_dmac_m_src_axi_wstrb
	wire          video_dmac_m_src_axi_wready;                                            // mm_interconnect_3:video_dmac_m_src_axi_wready -> video_dmac:m_src_axi_wready
	wire          video_dmac_m_src_axi_rid;                                               // mm_interconnect_3:video_dmac_m_src_axi_rid -> video_dmac:m_src_axi_rid
	wire          video_dmac_m_src_axi_rready;                                            // video_dmac:m_src_axi_rready -> mm_interconnect_3:video_dmac_m_src_axi_rready
	wire    [3:0] video_dmac_m_src_axi_awlen;                                             // video_dmac:m_src_axi_awlen -> mm_interconnect_3:video_dmac_m_src_axi_awlen
	wire          video_dmac_m_src_axi_wid;                                               // video_dmac:m_src_axi_wid -> mm_interconnect_3:video_dmac_m_src_axi_wid
	wire    [3:0] video_dmac_m_src_axi_arcache;                                           // video_dmac:m_src_axi_arcache -> mm_interconnect_3:video_dmac_m_src_axi_arcache
	wire          video_dmac_m_src_axi_wvalid;                                            // video_dmac:m_src_axi_wvalid -> mm_interconnect_3:video_dmac_m_src_axi_wvalid
	wire   [31:0] video_dmac_m_src_axi_araddr;                                            // video_dmac:m_src_axi_araddr -> mm_interconnect_3:video_dmac_m_src_axi_araddr
	wire    [2:0] video_dmac_m_src_axi_arprot;                                            // video_dmac:m_src_axi_arprot -> mm_interconnect_3:video_dmac_m_src_axi_arprot
	wire   [63:0] video_dmac_m_src_axi_wdata;                                             // video_dmac:m_src_axi_wdata -> mm_interconnect_3:video_dmac_m_src_axi_wdata
	wire          video_dmac_m_src_axi_arvalid;                                           // video_dmac:m_src_axi_arvalid -> mm_interconnect_3:video_dmac_m_src_axi_arvalid
	wire    [2:0] video_dmac_m_src_axi_awprot;                                            // video_dmac:m_src_axi_awprot -> mm_interconnect_3:video_dmac_m_src_axi_awprot
	wire    [3:0] video_dmac_m_src_axi_awcache;                                           // video_dmac:m_src_axi_awcache -> mm_interconnect_3:video_dmac_m_src_axi_awcache
	wire          video_dmac_m_src_axi_arid;                                              // video_dmac:m_src_axi_arid -> mm_interconnect_3:video_dmac_m_src_axi_arid
	wire    [1:0] video_dmac_m_src_axi_arlock;                                            // video_dmac:m_src_axi_arlock -> mm_interconnect_3:video_dmac_m_src_axi_arlock
	wire    [1:0] video_dmac_m_src_axi_awlock;                                            // video_dmac:m_src_axi_awlock -> mm_interconnect_3:video_dmac_m_src_axi_awlock
	wire   [31:0] video_dmac_m_src_axi_awaddr;                                            // video_dmac:m_src_axi_awaddr -> mm_interconnect_3:video_dmac_m_src_axi_awaddr
	wire    [1:0] video_dmac_m_src_axi_bresp;                                             // mm_interconnect_3:video_dmac_m_src_axi_bresp -> video_dmac:m_src_axi_bresp
	wire          video_dmac_m_src_axi_arready;                                           // mm_interconnect_3:video_dmac_m_src_axi_arready -> video_dmac:m_src_axi_arready
	wire   [63:0] video_dmac_m_src_axi_rdata;                                             // mm_interconnect_3:video_dmac_m_src_axi_rdata -> video_dmac:m_src_axi_rdata
	wire          video_dmac_m_src_axi_awready;                                           // mm_interconnect_3:video_dmac_m_src_axi_awready -> video_dmac:m_src_axi_awready
	wire    [1:0] video_dmac_m_src_axi_arburst;                                           // video_dmac:m_src_axi_arburst -> mm_interconnect_3:video_dmac_m_src_axi_arburst
	wire    [2:0] video_dmac_m_src_axi_arsize;                                            // video_dmac:m_src_axi_arsize -> mm_interconnect_3:video_dmac_m_src_axi_arsize
	wire          video_dmac_m_src_axi_bready;                                            // video_dmac:m_src_axi_bready -> mm_interconnect_3:video_dmac_m_src_axi_bready
	wire          video_dmac_m_src_axi_rlast;                                             // mm_interconnect_3:video_dmac_m_src_axi_rlast -> video_dmac:m_src_axi_rlast
	wire          video_dmac_m_src_axi_wlast;                                             // video_dmac:m_src_axi_wlast -> mm_interconnect_3:video_dmac_m_src_axi_wlast
	wire    [1:0] video_dmac_m_src_axi_rresp;                                             // mm_interconnect_3:video_dmac_m_src_axi_rresp -> video_dmac:m_src_axi_rresp
	wire          video_dmac_m_src_axi_awid;                                              // video_dmac:m_src_axi_awid -> mm_interconnect_3:video_dmac_m_src_axi_awid
	wire          video_dmac_m_src_axi_bid;                                               // mm_interconnect_3:video_dmac_m_src_axi_bid -> video_dmac:m_src_axi_bid
	wire          video_dmac_m_src_axi_bvalid;                                            // mm_interconnect_3:video_dmac_m_src_axi_bvalid -> video_dmac:m_src_axi_bvalid
	wire          video_dmac_m_src_axi_awvalid;                                           // video_dmac:m_src_axi_awvalid -> mm_interconnect_3:video_dmac_m_src_axi_awvalid
	wire          video_dmac_m_src_axi_rvalid;                                            // mm_interconnect_3:video_dmac_m_src_axi_rvalid -> video_dmac:m_src_axi_rvalid
	wire    [2:0] video_dmac_m_src_axi_awsize;                                            // video_dmac:m_src_axi_awsize -> mm_interconnect_3:video_dmac_m_src_axi_awsize
	wire    [1:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_awburst;                      // mm_interconnect_3:sys_hps_f2h_sdram0_data_awburst -> sys_hps:f2h_sdram0_AWBURST
	wire    [3:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_arlen;                        // mm_interconnect_3:sys_hps_f2h_sdram0_data_arlen -> sys_hps:f2h_sdram0_ARLEN
	wire    [7:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_wstrb;                        // mm_interconnect_3:sys_hps_f2h_sdram0_data_wstrb -> sys_hps:f2h_sdram0_WSTRB
	wire          mm_interconnect_3_sys_hps_f2h_sdram0_data_wready;                       // sys_hps:f2h_sdram0_WREADY -> mm_interconnect_3:sys_hps_f2h_sdram0_data_wready
	wire    [7:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_rid;                          // sys_hps:f2h_sdram0_RID -> mm_interconnect_3:sys_hps_f2h_sdram0_data_rid
	wire          mm_interconnect_3_sys_hps_f2h_sdram0_data_rready;                       // mm_interconnect_3:sys_hps_f2h_sdram0_data_rready -> sys_hps:f2h_sdram0_RREADY
	wire    [3:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_awlen;                        // mm_interconnect_3:sys_hps_f2h_sdram0_data_awlen -> sys_hps:f2h_sdram0_AWLEN
	wire    [7:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_wid;                          // mm_interconnect_3:sys_hps_f2h_sdram0_data_wid -> sys_hps:f2h_sdram0_WID
	wire    [3:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_arcache;                      // mm_interconnect_3:sys_hps_f2h_sdram0_data_arcache -> sys_hps:f2h_sdram0_ARCACHE
	wire          mm_interconnect_3_sys_hps_f2h_sdram0_data_wvalid;                       // mm_interconnect_3:sys_hps_f2h_sdram0_data_wvalid -> sys_hps:f2h_sdram0_WVALID
	wire   [31:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_araddr;                       // mm_interconnect_3:sys_hps_f2h_sdram0_data_araddr -> sys_hps:f2h_sdram0_ARADDR
	wire    [2:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_arprot;                       // mm_interconnect_3:sys_hps_f2h_sdram0_data_arprot -> sys_hps:f2h_sdram0_ARPROT
	wire    [2:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_awprot;                       // mm_interconnect_3:sys_hps_f2h_sdram0_data_awprot -> sys_hps:f2h_sdram0_AWPROT
	wire   [63:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_wdata;                        // mm_interconnect_3:sys_hps_f2h_sdram0_data_wdata -> sys_hps:f2h_sdram0_WDATA
	wire          mm_interconnect_3_sys_hps_f2h_sdram0_data_arvalid;                      // mm_interconnect_3:sys_hps_f2h_sdram0_data_arvalid -> sys_hps:f2h_sdram0_ARVALID
	wire    [3:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_awcache;                      // mm_interconnect_3:sys_hps_f2h_sdram0_data_awcache -> sys_hps:f2h_sdram0_AWCACHE
	wire    [7:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_arid;                         // mm_interconnect_3:sys_hps_f2h_sdram0_data_arid -> sys_hps:f2h_sdram0_ARID
	wire    [1:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_arlock;                       // mm_interconnect_3:sys_hps_f2h_sdram0_data_arlock -> sys_hps:f2h_sdram0_ARLOCK
	wire    [1:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_awlock;                       // mm_interconnect_3:sys_hps_f2h_sdram0_data_awlock -> sys_hps:f2h_sdram0_AWLOCK
	wire   [31:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_awaddr;                       // mm_interconnect_3:sys_hps_f2h_sdram0_data_awaddr -> sys_hps:f2h_sdram0_AWADDR
	wire    [1:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_bresp;                        // sys_hps:f2h_sdram0_BRESP -> mm_interconnect_3:sys_hps_f2h_sdram0_data_bresp
	wire          mm_interconnect_3_sys_hps_f2h_sdram0_data_arready;                      // sys_hps:f2h_sdram0_ARREADY -> mm_interconnect_3:sys_hps_f2h_sdram0_data_arready
	wire   [63:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_rdata;                        // sys_hps:f2h_sdram0_RDATA -> mm_interconnect_3:sys_hps_f2h_sdram0_data_rdata
	wire          mm_interconnect_3_sys_hps_f2h_sdram0_data_awready;                      // sys_hps:f2h_sdram0_AWREADY -> mm_interconnect_3:sys_hps_f2h_sdram0_data_awready
	wire    [1:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_arburst;                      // mm_interconnect_3:sys_hps_f2h_sdram0_data_arburst -> sys_hps:f2h_sdram0_ARBURST
	wire    [2:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_arsize;                       // mm_interconnect_3:sys_hps_f2h_sdram0_data_arsize -> sys_hps:f2h_sdram0_ARSIZE
	wire          mm_interconnect_3_sys_hps_f2h_sdram0_data_bready;                       // mm_interconnect_3:sys_hps_f2h_sdram0_data_bready -> sys_hps:f2h_sdram0_BREADY
	wire          mm_interconnect_3_sys_hps_f2h_sdram0_data_rlast;                        // sys_hps:f2h_sdram0_RLAST -> mm_interconnect_3:sys_hps_f2h_sdram0_data_rlast
	wire          mm_interconnect_3_sys_hps_f2h_sdram0_data_wlast;                        // mm_interconnect_3:sys_hps_f2h_sdram0_data_wlast -> sys_hps:f2h_sdram0_WLAST
	wire    [1:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_rresp;                        // sys_hps:f2h_sdram0_RRESP -> mm_interconnect_3:sys_hps_f2h_sdram0_data_rresp
	wire    [7:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_awid;                         // mm_interconnect_3:sys_hps_f2h_sdram0_data_awid -> sys_hps:f2h_sdram0_AWID
	wire    [7:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_bid;                          // sys_hps:f2h_sdram0_BID -> mm_interconnect_3:sys_hps_f2h_sdram0_data_bid
	wire          mm_interconnect_3_sys_hps_f2h_sdram0_data_bvalid;                       // sys_hps:f2h_sdram0_BVALID -> mm_interconnect_3:sys_hps_f2h_sdram0_data_bvalid
	wire    [2:0] mm_interconnect_3_sys_hps_f2h_sdram0_data_awsize;                       // mm_interconnect_3:sys_hps_f2h_sdram0_data_awsize -> sys_hps:f2h_sdram0_AWSIZE
	wire          mm_interconnect_3_sys_hps_f2h_sdram0_data_awvalid;                      // mm_interconnect_3:sys_hps_f2h_sdram0_data_awvalid -> sys_hps:f2h_sdram0_AWVALID
	wire          mm_interconnect_3_sys_hps_f2h_sdram0_data_rvalid;                       // sys_hps:f2h_sdram0_RVALID -> mm_interconnect_3:sys_hps_f2h_sdram0_data_rvalid
	wire          irq_mapper_receiver0_irq;                                               // video_dmac:irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                               // axi_adc_dma:irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                               // sys_gpio_bd:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                               // sys_spi:irq -> irq_mapper:receiver3_irq
	wire   [31:0] sys_hps_f2h_irq0_irq;                                                   // irq_mapper:sender_irq -> sys_hps:f2h_irq_p0
	wire   [31:0] sys_hps_f2h_irq1_irq;                                                   // irq_mapper_001:sender_irq -> sys_hps:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                                         // rst_controller:reset_out -> [adc_pwm_gen:s_axi_aresetn, axi_adc_dma:m_dest_axi_aresetn, axi_adc_dma:s_axi_aresetn, axi_ltc235x:s_axi_aresetn, axi_sysid_0:s_axi_aresetn, mm_interconnect_0:sys_int_mem_reset1_reset_bridge_in_reset_reset, mm_interconnect_1:sys_id_reset_reset_bridge_in_reset_reset, mm_interconnect_2:axi_adc_dma_m_dest_axi_reset_reset_bridge_in_reset_reset, pixel_clk_pll_reconfig:mgmt_reset, rst_translator:in_reset, sys_gpio_bd:reset_n, sys_gpio_in:reset_n, sys_gpio_out:reset_n, sys_id:reset_n, sys_int_mem:reset, sys_spi:reset_n, util_adc_pack:reset, vga_out:s_axi_aresetn, video_dmac:s_axi_aresetn]
	wire          rst_controller_reset_out_reset_req;                                     // rst_controller:reset_req -> [rst_translator:reset_req_in, sys_int_mem:reset_req]
	wire          rst_controller_001_reset_out_reset;                                     // rst_controller_001:reset_out -> [mm_interconnect_3:video_dmac_m_src_axi_reset_reset_bridge_in_reset_reset, video_dmac:m_src_axi_aresetn]
	wire          rst_controller_002_reset_out_reset;                                     // rst_controller_002:reset_out -> [mm_interconnect_0:sys_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sys_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_003_reset_out_reset;                                     // rst_controller_003:reset_out -> mm_interconnect_2:sys_hps_f2h_sdram1_data_agent_reset_sink_reset_bridge_in_reset_reset
	wire          rst_controller_004_reset_out_reset;                                     // rst_controller_004:reset_out -> mm_interconnect_3:video_dmac_m_src_axi_id_pad_clk_reset_reset_bridge_in_reset_reset

	axi_pwm_gen #(
		.ID             (0),
		.ASYNC_CLK_EN   (0),
		.N_PWMS         (1),
		.PWM_EXT_SYNC   (0),
		.EXT_ASYNC_SYNC (0),
		.PULSE_0_WIDTH  (1),
		.PULSE_1_WIDTH  (7),
		.PULSE_2_WIDTH  (7),
		.PULSE_3_WIDTH  (7),
		.PULSE_0_PERIOD (8),
		.PULSE_1_PERIOD (10),
		.PULSE_2_PERIOD (10),
		.PULSE_3_PERIOD (10),
		.PULSE_0_OFFSET (0),
		.PULSE_1_OFFSET (0),
		.PULSE_2_OFFSET (0),
		.PULSE_3_OFFSET (0)
	) adc_pwm_gen (
		.s_axi_aclk    (sys_clk_clk),                                 // s_axi_clock.clk
		.s_axi_aresetn (~rst_controller_reset_out_reset),             // s_axi_reset.reset_n
		.s_axi_awvalid (mm_interconnect_1_adc_pwm_gen_s_axi_awvalid), //       s_axi.awvalid
		.s_axi_awaddr  (mm_interconnect_1_adc_pwm_gen_s_axi_awaddr),  //            .awaddr
		.s_axi_awprot  (mm_interconnect_1_adc_pwm_gen_s_axi_awprot),  //            .awprot
		.s_axi_awready (mm_interconnect_1_adc_pwm_gen_s_axi_awready), //            .awready
		.s_axi_wvalid  (mm_interconnect_1_adc_pwm_gen_s_axi_wvalid),  //            .wvalid
		.s_axi_wdata   (mm_interconnect_1_adc_pwm_gen_s_axi_wdata),   //            .wdata
		.s_axi_wstrb   (mm_interconnect_1_adc_pwm_gen_s_axi_wstrb),   //            .wstrb
		.s_axi_wready  (mm_interconnect_1_adc_pwm_gen_s_axi_wready),  //            .wready
		.s_axi_bvalid  (mm_interconnect_1_adc_pwm_gen_s_axi_bvalid),  //            .bvalid
		.s_axi_bresp   (mm_interconnect_1_adc_pwm_gen_s_axi_bresp),   //            .bresp
		.s_axi_bready  (mm_interconnect_1_adc_pwm_gen_s_axi_bready),  //            .bready
		.s_axi_arvalid (mm_interconnect_1_adc_pwm_gen_s_axi_arvalid), //            .arvalid
		.s_axi_araddr  (mm_interconnect_1_adc_pwm_gen_s_axi_araddr),  //            .araddr
		.s_axi_arprot  (mm_interconnect_1_adc_pwm_gen_s_axi_arprot),  //            .arprot
		.s_axi_arready (mm_interconnect_1_adc_pwm_gen_s_axi_arready), //            .arready
		.s_axi_rvalid  (mm_interconnect_1_adc_pwm_gen_s_axi_rvalid),  //            .rvalid
		.s_axi_rresp   (mm_interconnect_1_adc_pwm_gen_s_axi_rresp),   //            .rresp
		.s_axi_rdata   (mm_interconnect_1_adc_pwm_gen_s_axi_rdata),   //            .rdata
		.s_axi_rready  (mm_interconnect_1_adc_pwm_gen_s_axi_rready),  //            .rready
		.ext_clk       (sys_clk_clk),                                 //  if_ext_clk.clk
		.ext_sync      (),                                            // if_ext_sync.ext_sync
		.pwm_0         (axi_ltc235x_cnv_if_pwm_0),                    //    if_pwm_0.pwm_0
		.pwm_1         (),                                            //    if_pwm_1.pwm_1
		.pwm_2         (),                                            //    if_pwm_2.pwm_2
		.pwm_3         ()                                             //    if_pwm_3.pwm_3
	);

	axi_dmac #(
		.ID                    (0),
		.DMA_LENGTH_WIDTH      (24),
		.FIFO_SIZE             (4),
		.MAX_BYTES_PER_BURST   (128),
		.DMA_TYPE_SRC          (2),
		.DMA_AXI_PROTOCOL_SRC  (1),
		.DMA_DATA_WIDTH_SRC    (256),
		.AXI_SLICE_SRC         (0),
		.DMA_TYPE_DEST         (0),
		.DMA_AXI_PROTOCOL_DEST (1),
		.DMA_DATA_WIDTH_DEST   (64),
		.AXI_SLICE_DEST        (0),
		.CYCLIC                (0),
		.DMA_2D_TRANSFER       (0),
		.SYNC_TRANSFER_START   (1),
		.ASYNC_CLK_REQ_SRC     (0),
		.ASYNC_CLK_SRC_DEST    (0),
		.ASYNC_CLK_DEST_REQ    (0),
		.ENABLE_DIAGNOSTICS_IF (0),
		.DMA_AXIS_ID_W         (8),
		.DMA_AXIS_DEST_W       (4)
	) axi_adc_dma (
		.s_axi_aclk             (sys_clk_clk),                                                                                                                                                                                                                                                           //         s_axi_clock.clk
		.s_axi_aresetn          (~rst_controller_reset_out_reset),                                                                                                                                                                                                                                       //         s_axi_reset.reset_n
		.s_axi_awvalid          (mm_interconnect_1_axi_adc_dma_s_axi_awvalid),                                                                                                                                                                                                                           //               s_axi.awvalid
		.s_axi_awaddr           (mm_interconnect_1_axi_adc_dma_s_axi_awaddr),                                                                                                                                                                                                                            //                    .awaddr
		.s_axi_awprot           (mm_interconnect_1_axi_adc_dma_s_axi_awprot),                                                                                                                                                                                                                            //                    .awprot
		.s_axi_awready          (mm_interconnect_1_axi_adc_dma_s_axi_awready),                                                                                                                                                                                                                           //                    .awready
		.s_axi_wvalid           (mm_interconnect_1_axi_adc_dma_s_axi_wvalid),                                                                                                                                                                                                                            //                    .wvalid
		.s_axi_wdata            (mm_interconnect_1_axi_adc_dma_s_axi_wdata),                                                                                                                                                                                                                             //                    .wdata
		.s_axi_wstrb            (mm_interconnect_1_axi_adc_dma_s_axi_wstrb),                                                                                                                                                                                                                             //                    .wstrb
		.s_axi_wready           (mm_interconnect_1_axi_adc_dma_s_axi_wready),                                                                                                                                                                                                                            //                    .wready
		.s_axi_bvalid           (mm_interconnect_1_axi_adc_dma_s_axi_bvalid),                                                                                                                                                                                                                            //                    .bvalid
		.s_axi_bresp            (mm_interconnect_1_axi_adc_dma_s_axi_bresp),                                                                                                                                                                                                                             //                    .bresp
		.s_axi_bready           (mm_interconnect_1_axi_adc_dma_s_axi_bready),                                                                                                                                                                                                                            //                    .bready
		.s_axi_arvalid          (mm_interconnect_1_axi_adc_dma_s_axi_arvalid),                                                                                                                                                                                                                           //                    .arvalid
		.s_axi_araddr           (mm_interconnect_1_axi_adc_dma_s_axi_araddr),                                                                                                                                                                                                                            //                    .araddr
		.s_axi_arprot           (mm_interconnect_1_axi_adc_dma_s_axi_arprot),                                                                                                                                                                                                                            //                    .arprot
		.s_axi_arready          (mm_interconnect_1_axi_adc_dma_s_axi_arready),                                                                                                                                                                                                                           //                    .arready
		.s_axi_rvalid           (mm_interconnect_1_axi_adc_dma_s_axi_rvalid),                                                                                                                                                                                                                            //                    .rvalid
		.s_axi_rresp            (mm_interconnect_1_axi_adc_dma_s_axi_rresp),                                                                                                                                                                                                                             //                    .rresp
		.s_axi_rdata            (mm_interconnect_1_axi_adc_dma_s_axi_rdata),                                                                                                                                                                                                                             //                    .rdata
		.s_axi_rready           (mm_interconnect_1_axi_adc_dma_s_axi_rready),                                                                                                                                                                                                                            //                    .rready
		.irq                    (irq_mapper_receiver1_irq),                                                                                                                                                                                                                                              //    interrupt_sender.irq
		.m_dest_axi_aclk        (sys_clk_clk),                                                                                                                                                                                                                                                           //    m_dest_axi_clock.clk
		.m_dest_axi_aresetn     (~rst_controller_reset_out_reset),                                                                                                                                                                                                                                       //    m_dest_axi_reset.reset_n
		.fifo_wr_clk            (sys_clk_clk),                                                                                                                                                                                                                                                           //      if_fifo_wr_clk.clk
		.fifo_wr_en             (util_adc_pack_if_packed_fifo_wr_en_valid),                                                                                                                                                                                                                              //       if_fifo_wr_en.valid
		.fifo_wr_din            (util_adc_pack_if_packed_fifo_wr_data_data),                                                                                                                                                                                                                             //      if_fifo_wr_din.data
		.fifo_wr_overflow       (axi_adc_dma_if_fifo_wr_overflow_ovf),                                                                                                                                                                                                                                   // if_fifo_wr_overflow.ovf
		.fifo_wr_sync           (util_adc_pack_if_packed_fifo_wr_sync_sync),                                                                                                                                                                                                                             //     if_fifo_wr_sync.sync
		.fifo_wr_xfer_req       (),                                                                                                                                                                                                                                                                      // if_fifo_wr_xfer_req.xfer_req
		.m_dest_axi_awvalid     (axi_adc_dma_m_dest_axi_awvalid),                                                                                                                                                                                                                                        //          m_dest_axi.awvalid
		.m_dest_axi_awaddr      (axi_adc_dma_m_dest_axi_awaddr),                                                                                                                                                                                                                                         //                    .awaddr
		.m_dest_axi_awready     (axi_adc_dma_m_dest_axi_awready),                                                                                                                                                                                                                                        //                    .awready
		.m_dest_axi_wvalid      (axi_adc_dma_m_dest_axi_wvalid),                                                                                                                                                                                                                                         //                    .wvalid
		.m_dest_axi_wdata       (axi_adc_dma_m_dest_axi_wdata),                                                                                                                                                                                                                                          //                    .wdata
		.m_dest_axi_wstrb       (axi_adc_dma_m_dest_axi_wstrb),                                                                                                                                                                                                                                          //                    .wstrb
		.m_dest_axi_wready      (axi_adc_dma_m_dest_axi_wready),                                                                                                                                                                                                                                         //                    .wready
		.m_dest_axi_bvalid      (axi_adc_dma_m_dest_axi_bvalid),                                                                                                                                                                                                                                         //                    .bvalid
		.m_dest_axi_bresp       (axi_adc_dma_m_dest_axi_bresp),                                                                                                                                                                                                                                          //                    .bresp
		.m_dest_axi_bready      (axi_adc_dma_m_dest_axi_bready),                                                                                                                                                                                                                                         //                    .bready
		.m_dest_axi_arvalid     (axi_adc_dma_m_dest_axi_arvalid),                                                                                                                                                                                                                                        //                    .arvalid
		.m_dest_axi_araddr      (axi_adc_dma_m_dest_axi_araddr),                                                                                                                                                                                                                                         //                    .araddr
		.m_dest_axi_arready     (axi_adc_dma_m_dest_axi_arready),                                                                                                                                                                                                                                        //                    .arready
		.m_dest_axi_rvalid      (axi_adc_dma_m_dest_axi_rvalid),                                                                                                                                                                                                                                         //                    .rvalid
		.m_dest_axi_rresp       (axi_adc_dma_m_dest_axi_rresp),                                                                                                                                                                                                                                          //                    .rresp
		.m_dest_axi_rdata       (axi_adc_dma_m_dest_axi_rdata),                                                                                                                                                                                                                                          //                    .rdata
		.m_dest_axi_rready      (axi_adc_dma_m_dest_axi_rready),                                                                                                                                                                                                                                         //                    .rready
		.m_dest_axi_awlen       (axi_adc_dma_m_dest_axi_awlen),                                                                                                                                                                                                                                          //                    .awlen
		.m_dest_axi_awsize      (axi_adc_dma_m_dest_axi_awsize),                                                                                                                                                                                                                                         //                    .awsize
		.m_dest_axi_awburst     (axi_adc_dma_m_dest_axi_awburst),                                                                                                                                                                                                                                        //                    .awburst
		.m_dest_axi_awcache     (axi_adc_dma_m_dest_axi_awcache),                                                                                                                                                                                                                                        //                    .awcache
		.m_dest_axi_awprot      (axi_adc_dma_m_dest_axi_awprot),                                                                                                                                                                                                                                         //                    .awprot
		.m_dest_axi_wlast       (axi_adc_dma_m_dest_axi_wlast),                                                                                                                                                                                                                                          //                    .wlast
		.m_dest_axi_arlen       (axi_adc_dma_m_dest_axi_arlen),                                                                                                                                                                                                                                          //                    .arlen
		.m_dest_axi_arsize      (axi_adc_dma_m_dest_axi_arsize),                                                                                                                                                                                                                                         //                    .arsize
		.m_dest_axi_arburst     (axi_adc_dma_m_dest_axi_arburst),                                                                                                                                                                                                                                        //                    .arburst
		.m_dest_axi_arcache     (axi_adc_dma_m_dest_axi_arcache),                                                                                                                                                                                                                                        //                    .arcache
		.m_dest_axi_arprot      (axi_adc_dma_m_dest_axi_arprot),                                                                                                                                                                                                                                         //                    .arprot
		.m_dest_axi_awid        (axi_adc_dma_m_dest_axi_awid),                                                                                                                                                                                                                                           //                    .awid
		.m_dest_axi_awlock      (axi_adc_dma_m_dest_axi_awlock),                                                                                                                                                                                                                                         //                    .awlock
		.m_dest_axi_wid         (axi_adc_dma_m_dest_axi_wid),                                                                                                                                                                                                                                            //                    .wid
		.m_dest_axi_arid        (axi_adc_dma_m_dest_axi_arid),                                                                                                                                                                                                                                           //                    .arid
		.m_dest_axi_arlock      (axi_adc_dma_m_dest_axi_arlock),                                                                                                                                                                                                                                         //                    .arlock
		.m_dest_axi_rid         (axi_adc_dma_m_dest_axi_rid),                                                                                                                                                                                                                                            //                    .rid
		.m_dest_axi_bid         (axi_adc_dma_m_dest_axi_bid),                                                                                                                                                                                                                                            //                    .bid
		.m_dest_axi_rlast       (axi_adc_dma_m_dest_axi_rlast),                                                                                                                                                                                                                                          //                    .rlast
		.m_src_axi_aclk         (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.m_src_axi_aresetn      (1'b1),                                                                                                                                                                                                                                                                  //         (terminated)
		.m_axis_aclk            (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.m_axis_xfer_req        (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_axis_valid           (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_axis_last            (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_axis_ready           (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.m_axis_data            (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_axis_user            (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_axis_id              (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_axis_dest            (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_axis_strb            (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_axis_keep            (),                                                                                                                                                                                                                                                                      //         (terminated)
		.s_axis_aclk            (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.s_axis_xfer_req        (),                                                                                                                                                                                                                                                                      //         (terminated)
		.s_axis_valid           (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.s_axis_last            (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.s_axis_ready           (),                                                                                                                                                                                                                                                                      //         (terminated)
		.s_axis_data            (256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //         (terminated)
		.s_axis_user            (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.s_axis_id              (8'b00000000),                                                                                                                                                                                                                                                           //         (terminated)
		.s_axis_dest            (4'b0000),                                                                                                                                                                                                                                                               //         (terminated)
		.s_axis_strb            (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  //         (terminated)
		.s_axis_keep            (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  //         (terminated)
		.fifo_rd_clk            (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.fifo_rd_en             (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.fifo_rd_valid          (),                                                                                                                                                                                                                                                                      //         (terminated)
		.fifo_rd_dout           (),                                                                                                                                                                                                                                                                      //         (terminated)
		.fifo_rd_underflow      (),                                                                                                                                                                                                                                                                      //         (terminated)
		.fifo_rd_xfer_req       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.dest_diag_level_bursts (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_awvalid      (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_awaddr       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_awready      (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.m_src_axi_wvalid       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_wdata        (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_wstrb        (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_wready       (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.m_src_axi_bvalid       (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.m_src_axi_bresp        (2'b00),                                                                                                                                                                                                                                                                 //         (terminated)
		.m_src_axi_bready       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_arvalid      (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_araddr       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_arready      (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.m_src_axi_rvalid       (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.m_src_axi_rresp        (2'b00),                                                                                                                                                                                                                                                                 //         (terminated)
		.m_src_axi_rdata        (256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //         (terminated)
		.m_src_axi_rready       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_awlen        (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_awsize       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_awburst      (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_awcache      (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_awprot       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_wlast        (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_arlen        (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_arsize       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_arburst      (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_arcache      (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_arprot       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_awid         (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_awlock       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_wid          (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_arid         (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_arlock       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.m_src_axi_rid          (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.m_src_axi_bid          (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.m_src_axi_rlast        (1'b0)                                                                                                                                                                                                                                                                   //         (terminated)
	);

	axi_ltc235x #(
		.ID              (0),
		.LVDS_CMOS_N     (0),
		.LANE_0_ENABLE   (1),
		.LANE_1_ENABLE   (1),
		.LANE_2_ENABLE   (1),
		.LANE_3_ENABLE   (1),
		.LANE_4_ENABLE   (1),
		.LANE_5_ENABLE   (1),
		.LANE_6_ENABLE   (1),
		.LANE_7_ENABLE   (1),
		.NUM_CHANNELS    (8),
		.DATA_WIDTH      (18),
		.SOFTSPAN_NEXT   (16777215),
		.EXTERNAL_CLK    (0),
		.FPGA_TECHNOLOGY (101),
		.FPGA_FAMILY     (1),
		.SPEED_GRADE     (8),
		.DEV_PACKAGE     (3)
	) axi_ltc235x (
		.busy          (axi_ltc235x_device_if_busy),                  //       device_if.busy
		.lvds_cmos_n   (axi_ltc235x_device_if_lvds_cmos_n),           //                .lvds_cmos_n
		.cs_n          (axi_ltc235x_device_if_cs_n),                  //                .cs_n
		.pd            (axi_ltc235x_device_if_pd),                    //                .pd
		.scki          (axi_ltc235x_device_if_scki),                  //                .scki
		.scko          (axi_ltc235x_device_if_scko),                  //                .scko
		.sdi           (axi_ltc235x_device_if_sdi),                   //                .sdi
		.sdo_0         (axi_ltc235x_device_if_sdo_0),                 //                .sdo_0
		.sdo_1         (axi_ltc235x_device_if_sdo_1),                 //                .sdo_1
		.sdo_2         (axi_ltc235x_device_if_sdo_2),                 //                .sdo_2
		.sdo_3         (axi_ltc235x_device_if_sdo_3),                 //                .sdo_3
		.sdo_4         (axi_ltc235x_device_if_sdo_4),                 //                .sdo_4
		.sdo_5         (axi_ltc235x_device_if_sdo_5),                 //                .sdo_5
		.sdo_6         (axi_ltc235x_device_if_sdo_6),                 //                .sdo_6
		.sdo_7         (axi_ltc235x_device_if_sdo_7),                 //                .sdo_7
		.external_clk  (sys_clk_clk),                                 // if_external_clk.clk
		.s_axi_aclk    (sys_clk_clk),                                 //     s_axi_clock.clk
		.s_axi_aresetn (~rst_controller_reset_out_reset),             //     s_axi_reset.reset_n
		.s_axi_awvalid (mm_interconnect_1_axi_ltc235x_s_axi_awvalid), //           s_axi.awvalid
		.s_axi_awaddr  (mm_interconnect_1_axi_ltc235x_s_axi_awaddr),  //                .awaddr
		.s_axi_awprot  (mm_interconnect_1_axi_ltc235x_s_axi_awprot),  //                .awprot
		.s_axi_awready (mm_interconnect_1_axi_ltc235x_s_axi_awready), //                .awready
		.s_axi_wvalid  (mm_interconnect_1_axi_ltc235x_s_axi_wvalid),  //                .wvalid
		.s_axi_wdata   (mm_interconnect_1_axi_ltc235x_s_axi_wdata),   //                .wdata
		.s_axi_wstrb   (mm_interconnect_1_axi_ltc235x_s_axi_wstrb),   //                .wstrb
		.s_axi_wready  (mm_interconnect_1_axi_ltc235x_s_axi_wready),  //                .wready
		.s_axi_bvalid  (mm_interconnect_1_axi_ltc235x_s_axi_bvalid),  //                .bvalid
		.s_axi_bresp   (mm_interconnect_1_axi_ltc235x_s_axi_bresp),   //                .bresp
		.s_axi_bready  (mm_interconnect_1_axi_ltc235x_s_axi_bready),  //                .bready
		.s_axi_arvalid (mm_interconnect_1_axi_ltc235x_s_axi_arvalid), //                .arvalid
		.s_axi_araddr  (mm_interconnect_1_axi_ltc235x_s_axi_araddr),  //                .araddr
		.s_axi_arprot  (mm_interconnect_1_axi_ltc235x_s_axi_arprot),  //                .arprot
		.s_axi_arready (mm_interconnect_1_axi_ltc235x_s_axi_arready), //                .arready
		.s_axi_rvalid  (mm_interconnect_1_axi_ltc235x_s_axi_rvalid),  //                .rvalid
		.s_axi_rresp   (mm_interconnect_1_axi_ltc235x_s_axi_rresp),   //                .rresp
		.s_axi_rdata   (mm_interconnect_1_axi_ltc235x_s_axi_rdata),   //                .rdata
		.s_axi_rready  (mm_interconnect_1_axi_ltc235x_s_axi_rready),  //                .rready
		.adc_dovf      (util_adc_pack_if_fifo_wr_overflow_ovf),       //     if_adc_dovf.ovf
		.adc_enable_0  (axi_ltc235x_adc_ch_0_enable),                 //        adc_ch_0.enable
		.adc_valid_0   (axi_ltc235x_adc_ch_0_valid),                  //                .valid
		.adc_data_0    (axi_ltc235x_adc_ch_0_data),                   //                .data
		.adc_enable_1  (axi_ltc235x_adc_ch_1_enable),                 //        adc_ch_1.enable
		.adc_valid_1   (axi_ltc235x_adc_ch_1_valid),                  //                .valid
		.adc_data_1    (axi_ltc235x_adc_ch_1_data),                   //                .data
		.adc_enable_2  (axi_ltc235x_adc_ch_2_enable),                 //        adc_ch_2.enable
		.adc_valid_2   (axi_ltc235x_adc_ch_2_valid),                  //                .valid
		.adc_data_2    (axi_ltc235x_adc_ch_2_data),                   //                .data
		.adc_enable_3  (axi_ltc235x_adc_ch_3_enable),                 //        adc_ch_3.enable
		.adc_valid_3   (axi_ltc235x_adc_ch_3_valid),                  //                .valid
		.adc_data_3    (axi_ltc235x_adc_ch_3_data),                   //                .data
		.adc_enable_4  (axi_ltc235x_adc_ch_4_enable),                 //        adc_ch_4.enable
		.adc_valid_4   (axi_ltc235x_adc_ch_4_valid),                  //                .valid
		.adc_data_4    (axi_ltc235x_adc_ch_4_data),                   //                .data
		.adc_enable_5  (axi_ltc235x_adc_ch_5_enable),                 //        adc_ch_5.enable
		.adc_valid_5   (axi_ltc235x_adc_ch_5_valid),                  //                .valid
		.adc_data_5    (axi_ltc235x_adc_ch_5_data),                   //                .data
		.adc_enable_6  (axi_ltc235x_adc_ch_6_enable),                 //        adc_ch_6.enable
		.adc_valid_6   (axi_ltc235x_adc_ch_6_valid),                  //                .valid
		.adc_data_6    (axi_ltc235x_adc_ch_6_data),                   //                .data
		.adc_enable_7  (axi_ltc235x_adc_ch_7_enable),                 //        adc_ch_7.enable
		.adc_valid_7   (axi_ltc235x_adc_ch_7_valid),                  //                .valid
		.adc_data_7    (axi_ltc235x_adc_ch_7_data)                    //                .data
	);

	axi_sysid #(
		.ROM_WIDTH     (32),
		.ROM_ADDR_BITS (9)
	) axi_sysid_0 (
		.s_axi_aclk    (sys_clk_clk),                                 //     s_axi_clock.clk
		.s_axi_aresetn (~rst_controller_reset_out_reset),             //     s_axi_reset.reset_n
		.s_axi_awvalid (mm_interconnect_1_axi_sysid_0_s_axi_awvalid), //           s_axi.awvalid
		.s_axi_awaddr  (mm_interconnect_1_axi_sysid_0_s_axi_awaddr),  //                .awaddr
		.s_axi_awprot  (mm_interconnect_1_axi_sysid_0_s_axi_awprot),  //                .awprot
		.s_axi_awready (mm_interconnect_1_axi_sysid_0_s_axi_awready), //                .awready
		.s_axi_wvalid  (mm_interconnect_1_axi_sysid_0_s_axi_wvalid),  //                .wvalid
		.s_axi_wdata   (mm_interconnect_1_axi_sysid_0_s_axi_wdata),   //                .wdata
		.s_axi_wstrb   (mm_interconnect_1_axi_sysid_0_s_axi_wstrb),   //                .wstrb
		.s_axi_wready  (mm_interconnect_1_axi_sysid_0_s_axi_wready),  //                .wready
		.s_axi_bvalid  (mm_interconnect_1_axi_sysid_0_s_axi_bvalid),  //                .bvalid
		.s_axi_bresp   (mm_interconnect_1_axi_sysid_0_s_axi_bresp),   //                .bresp
		.s_axi_bready  (mm_interconnect_1_axi_sysid_0_s_axi_bready),  //                .bready
		.s_axi_arvalid (mm_interconnect_1_axi_sysid_0_s_axi_arvalid), //                .arvalid
		.s_axi_araddr  (mm_interconnect_1_axi_sysid_0_s_axi_araddr),  //                .araddr
		.s_axi_arprot  (mm_interconnect_1_axi_sysid_0_s_axi_arprot),  //                .arprot
		.s_axi_arready (mm_interconnect_1_axi_sysid_0_s_axi_arready), //                .arready
		.s_axi_rvalid  (mm_interconnect_1_axi_sysid_0_s_axi_rvalid),  //                .rvalid
		.s_axi_rresp   (mm_interconnect_1_axi_sysid_0_s_axi_rresp),   //                .rresp
		.s_axi_rdata   (mm_interconnect_1_axi_sysid_0_s_axi_rdata),   //                .rdata
		.s_axi_rready  (mm_interconnect_1_axi_sysid_0_s_axi_rready),  //                .rready
		.sys_rom_data  (rom_sys_0_if_rom_data_rom_data),              // if_sys_rom_data.rom_data
		.pr_rom_data   (pr_rom_data_nc_rom_data),                     //  if_pr_rom_data.rom_data
		.rom_addr      (axi_sysid_0_if_rom_addr_rom_addr)             //     if_rom_addr.rom_addr
	);

	system_bd_pixel_clk_pll pixel_clk_pll (
		.refclk            (sys_clk_clk),                                            //            refclk.clk
		.rst               (~sys_rst_reset_n),                                       //             reset.reset
		.outclk_0          (pixel_clk_pll_outclk0_clk),                              //           outclk0.clk
		.outclk_1          (pixel_clk_pll_outclk1_clk),                              //           outclk1.clk
		.reconfig_to_pll   (pixel_clk_pll_reconfig_reconfig_to_pll_reconfig_to_pll), //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pixel_clk_pll_reconfig_from_pll_reconfig_from_pll),      // reconfig_from_pll.reconfig_from_pll
		.locked            ()                                                        //       (terminated)
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) pixel_clk_pll_reconfig (
		.mgmt_clk          (sys_clk_clk),                                                            //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_reset_out_reset),                                         //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (pixel_clk_pll_reconfig_reconfig_to_pll_reconfig_to_pll),                 //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pixel_clk_pll_reconfig_from_pll_reconfig_from_pll),                      // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                                 //       (terminated)
	);

	sysid_rom #(
		.ROM_WIDTH     (32),
		.ROM_ADDR_BITS (9),
		.PATH_TO_FILE  ("/home/guest/jemfgeronimo_workspace/ltc235x_hw_test/projects/dc2677a/c5soc/mem_init_sys.txt")
	) rom_sys_0 (
		.clk      (sys_clk_clk),                      //      if_clk.clk
		.rom_data (rom_sys_0_if_rom_data_rom_data),   // if_rom_data.rom_data
		.rom_addr (axi_sysid_0_if_rom_addr_rom_addr)  // if_rom_addr.rom_addr
	);

	system_bd_sys_gpio_bd sys_gpio_bd (
		.clk        (sys_clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_sys_gpio_bd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sys_gpio_bd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sys_gpio_bd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sys_gpio_bd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sys_gpio_bd_s1_readdata),   //                    .readdata
		.in_port    (sys_gpio_bd_in_port),                         // external_connection.export
		.out_port   (sys_gpio_bd_out_port),                        //                    .export
		.irq        (irq_mapper_receiver2_irq)                     //                 irq.irq
	);

	system_bd_sys_gpio_in sys_gpio_in (
		.clk        (sys_clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_sys_gpio_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sys_gpio_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sys_gpio_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sys_gpio_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sys_gpio_in_s1_readdata),   //                    .readdata
		.in_port    (sys_gpio_in_export),                          // external_connection.export
		.irq        ()                                             //                 irq.irq
	);

	system_bd_sys_gpio_out sys_gpio_out (
		.clk        (sys_clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_1_sys_gpio_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sys_gpio_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sys_gpio_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sys_gpio_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sys_gpio_out_s1_readdata),   //                    .readdata
		.out_port   (sys_gpio_out_export)                           // external_connection.export
	);

	system_bd_sys_hps #(
		.F2S_Width (2),
		.S2F_Width (2)
	) sys_hps (
		.h2f_user0_clk            (sys_hps_h2f_user0_clock_clk),                       //   h2f_user0_clock.clk
		.i2c0_scl                 (sys_hps_i2c0_scl_in_clk),                           //       i2c0_scl_in.clk
		.i2c0_out_clk             (sys_hps_i2c0_clk_clk),                              //          i2c0_clk.clk
		.i2c0_out_data            (sys_hps_i2c0_out_data),                             //              i2c0.out_data
		.i2c0_sda                 (sys_hps_i2c0_sda),                                  //                  .sda
		.mem_a                    (sys_hps_memory_mem_a),                              //            memory.mem_a
		.mem_ba                   (sys_hps_memory_mem_ba),                             //                  .mem_ba
		.mem_ck                   (sys_hps_memory_mem_ck),                             //                  .mem_ck
		.mem_ck_n                 (sys_hps_memory_mem_ck_n),                           //                  .mem_ck_n
		.mem_cke                  (sys_hps_memory_mem_cke),                            //                  .mem_cke
		.mem_cs_n                 (sys_hps_memory_mem_cs_n),                           //                  .mem_cs_n
		.mem_ras_n                (sys_hps_memory_mem_ras_n),                          //                  .mem_ras_n
		.mem_cas_n                (sys_hps_memory_mem_cas_n),                          //                  .mem_cas_n
		.mem_we_n                 (sys_hps_memory_mem_we_n),                           //                  .mem_we_n
		.mem_reset_n              (sys_hps_memory_mem_reset_n),                        //                  .mem_reset_n
		.mem_dq                   (sys_hps_memory_mem_dq),                             //                  .mem_dq
		.mem_dqs                  (sys_hps_memory_mem_dqs),                            //                  .mem_dqs
		.mem_dqs_n                (sys_hps_memory_mem_dqs_n),                          //                  .mem_dqs_n
		.mem_odt                  (sys_hps_memory_mem_odt),                            //                  .mem_odt
		.mem_dm                   (sys_hps_memory_mem_dm),                             //                  .mem_dm
		.oct_rzqin                (sys_hps_memory_oct_rzqin),                          //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (sys_hps_hps_io_hps_io_emac1_inst_TX_CLK),           //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (sys_hps_hps_io_hps_io_emac1_inst_TXD0),             //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (sys_hps_hps_io_hps_io_emac1_inst_TXD1),             //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (sys_hps_hps_io_hps_io_emac1_inst_TXD2),             //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (sys_hps_hps_io_hps_io_emac1_inst_TXD3),             //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (sys_hps_hps_io_hps_io_emac1_inst_RXD0),             //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (sys_hps_hps_io_hps_io_emac1_inst_MDIO),             //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (sys_hps_hps_io_hps_io_emac1_inst_MDC),              //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (sys_hps_hps_io_hps_io_emac1_inst_RX_CTL),           //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (sys_hps_hps_io_hps_io_emac1_inst_TX_CTL),           //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (sys_hps_hps_io_hps_io_emac1_inst_RX_CLK),           //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (sys_hps_hps_io_hps_io_emac1_inst_RXD1),             //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (sys_hps_hps_io_hps_io_emac1_inst_RXD2),             //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (sys_hps_hps_io_hps_io_emac1_inst_RXD3),             //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (sys_hps_hps_io_hps_io_qspi_inst_IO0),               //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (sys_hps_hps_io_hps_io_qspi_inst_IO1),               //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (sys_hps_hps_io_hps_io_qspi_inst_IO2),               //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (sys_hps_hps_io_hps_io_qspi_inst_IO3),               //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (sys_hps_hps_io_hps_io_qspi_inst_SS0),               //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (sys_hps_hps_io_hps_io_qspi_inst_CLK),               //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (sys_hps_hps_io_hps_io_sdio_inst_CMD),               //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (sys_hps_hps_io_hps_io_sdio_inst_D0),                //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (sys_hps_hps_io_hps_io_sdio_inst_D1),                //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (sys_hps_hps_io_hps_io_sdio_inst_CLK),               //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (sys_hps_hps_io_hps_io_sdio_inst_D2),                //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (sys_hps_hps_io_hps_io_sdio_inst_D3),                //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (sys_hps_hps_io_hps_io_usb1_inst_D0),                //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (sys_hps_hps_io_hps_io_usb1_inst_D1),                //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (sys_hps_hps_io_hps_io_usb1_inst_D2),                //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (sys_hps_hps_io_hps_io_usb1_inst_D3),                //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (sys_hps_hps_io_hps_io_usb1_inst_D4),                //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (sys_hps_hps_io_hps_io_usb1_inst_D5),                //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (sys_hps_hps_io_hps_io_usb1_inst_D6),                //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (sys_hps_hps_io_hps_io_usb1_inst_D7),                //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (sys_hps_hps_io_hps_io_usb1_inst_CLK),               //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (sys_hps_hps_io_hps_io_usb1_inst_STP),               //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (sys_hps_hps_io_hps_io_usb1_inst_DIR),               //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (sys_hps_hps_io_hps_io_usb1_inst_NXT),               //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (sys_hps_hps_io_hps_io_spim1_inst_CLK),              //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (sys_hps_hps_io_hps_io_spim1_inst_MOSI),             //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (sys_hps_hps_io_hps_io_spim1_inst_MISO),             //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (sys_hps_hps_io_hps_io_spim1_inst_SS0),              //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (sys_hps_hps_io_hps_io_uart0_inst_RX),               //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (sys_hps_hps_io_hps_io_uart0_inst_TX),               //                  .hps_io_uart0_inst_TX
		.h2f_rst_n                (sys_hps_h2f_reset_reset_n),                         //         h2f_reset.reset_n
		.f2h_sdram0_clk           (pixel_clk_pll_outclk1_clk),                         //  f2h_sdram0_clock.clk
		.f2h_sdram0_ARADDR        (mm_interconnect_3_sys_hps_f2h_sdram0_data_araddr),  //   f2h_sdram0_data.araddr
		.f2h_sdram0_ARLEN         (mm_interconnect_3_sys_hps_f2h_sdram0_data_arlen),   //                  .arlen
		.f2h_sdram0_ARID          (mm_interconnect_3_sys_hps_f2h_sdram0_data_arid),    //                  .arid
		.f2h_sdram0_ARSIZE        (mm_interconnect_3_sys_hps_f2h_sdram0_data_arsize),  //                  .arsize
		.f2h_sdram0_ARBURST       (mm_interconnect_3_sys_hps_f2h_sdram0_data_arburst), //                  .arburst
		.f2h_sdram0_ARLOCK        (mm_interconnect_3_sys_hps_f2h_sdram0_data_arlock),  //                  .arlock
		.f2h_sdram0_ARPROT        (mm_interconnect_3_sys_hps_f2h_sdram0_data_arprot),  //                  .arprot
		.f2h_sdram0_ARVALID       (mm_interconnect_3_sys_hps_f2h_sdram0_data_arvalid), //                  .arvalid
		.f2h_sdram0_ARCACHE       (mm_interconnect_3_sys_hps_f2h_sdram0_data_arcache), //                  .arcache
		.f2h_sdram0_AWADDR        (mm_interconnect_3_sys_hps_f2h_sdram0_data_awaddr),  //                  .awaddr
		.f2h_sdram0_AWLEN         (mm_interconnect_3_sys_hps_f2h_sdram0_data_awlen),   //                  .awlen
		.f2h_sdram0_AWID          (mm_interconnect_3_sys_hps_f2h_sdram0_data_awid),    //                  .awid
		.f2h_sdram0_AWSIZE        (mm_interconnect_3_sys_hps_f2h_sdram0_data_awsize),  //                  .awsize
		.f2h_sdram0_AWBURST       (mm_interconnect_3_sys_hps_f2h_sdram0_data_awburst), //                  .awburst
		.f2h_sdram0_AWLOCK        (mm_interconnect_3_sys_hps_f2h_sdram0_data_awlock),  //                  .awlock
		.f2h_sdram0_AWPROT        (mm_interconnect_3_sys_hps_f2h_sdram0_data_awprot),  //                  .awprot
		.f2h_sdram0_AWVALID       (mm_interconnect_3_sys_hps_f2h_sdram0_data_awvalid), //                  .awvalid
		.f2h_sdram0_AWCACHE       (mm_interconnect_3_sys_hps_f2h_sdram0_data_awcache), //                  .awcache
		.f2h_sdram0_BRESP         (mm_interconnect_3_sys_hps_f2h_sdram0_data_bresp),   //                  .bresp
		.f2h_sdram0_BID           (mm_interconnect_3_sys_hps_f2h_sdram0_data_bid),     //                  .bid
		.f2h_sdram0_BVALID        (mm_interconnect_3_sys_hps_f2h_sdram0_data_bvalid),  //                  .bvalid
		.f2h_sdram0_BREADY        (mm_interconnect_3_sys_hps_f2h_sdram0_data_bready),  //                  .bready
		.f2h_sdram0_ARREADY       (mm_interconnect_3_sys_hps_f2h_sdram0_data_arready), //                  .arready
		.f2h_sdram0_AWREADY       (mm_interconnect_3_sys_hps_f2h_sdram0_data_awready), //                  .awready
		.f2h_sdram0_RREADY        (mm_interconnect_3_sys_hps_f2h_sdram0_data_rready),  //                  .rready
		.f2h_sdram0_RDATA         (mm_interconnect_3_sys_hps_f2h_sdram0_data_rdata),   //                  .rdata
		.f2h_sdram0_RRESP         (mm_interconnect_3_sys_hps_f2h_sdram0_data_rresp),   //                  .rresp
		.f2h_sdram0_RLAST         (mm_interconnect_3_sys_hps_f2h_sdram0_data_rlast),   //                  .rlast
		.f2h_sdram0_RID           (mm_interconnect_3_sys_hps_f2h_sdram0_data_rid),     //                  .rid
		.f2h_sdram0_RVALID        (mm_interconnect_3_sys_hps_f2h_sdram0_data_rvalid),  //                  .rvalid
		.f2h_sdram0_WLAST         (mm_interconnect_3_sys_hps_f2h_sdram0_data_wlast),   //                  .wlast
		.f2h_sdram0_WVALID        (mm_interconnect_3_sys_hps_f2h_sdram0_data_wvalid),  //                  .wvalid
		.f2h_sdram0_WDATA         (mm_interconnect_3_sys_hps_f2h_sdram0_data_wdata),   //                  .wdata
		.f2h_sdram0_WSTRB         (mm_interconnect_3_sys_hps_f2h_sdram0_data_wstrb),   //                  .wstrb
		.f2h_sdram0_WREADY        (mm_interconnect_3_sys_hps_f2h_sdram0_data_wready),  //                  .wready
		.f2h_sdram0_WID           (mm_interconnect_3_sys_hps_f2h_sdram0_data_wid),     //                  .wid
		.f2h_sdram1_clk           (sys_hps_h2f_user0_clock_clk),                       //  f2h_sdram1_clock.clk
		.f2h_sdram1_ARADDR        (mm_interconnect_2_sys_hps_f2h_sdram1_data_araddr),  //   f2h_sdram1_data.araddr
		.f2h_sdram1_ARLEN         (mm_interconnect_2_sys_hps_f2h_sdram1_data_arlen),   //                  .arlen
		.f2h_sdram1_ARID          (mm_interconnect_2_sys_hps_f2h_sdram1_data_arid),    //                  .arid
		.f2h_sdram1_ARSIZE        (mm_interconnect_2_sys_hps_f2h_sdram1_data_arsize),  //                  .arsize
		.f2h_sdram1_ARBURST       (mm_interconnect_2_sys_hps_f2h_sdram1_data_arburst), //                  .arburst
		.f2h_sdram1_ARLOCK        (mm_interconnect_2_sys_hps_f2h_sdram1_data_arlock),  //                  .arlock
		.f2h_sdram1_ARPROT        (mm_interconnect_2_sys_hps_f2h_sdram1_data_arprot),  //                  .arprot
		.f2h_sdram1_ARVALID       (mm_interconnect_2_sys_hps_f2h_sdram1_data_arvalid), //                  .arvalid
		.f2h_sdram1_ARCACHE       (mm_interconnect_2_sys_hps_f2h_sdram1_data_arcache), //                  .arcache
		.f2h_sdram1_AWADDR        (mm_interconnect_2_sys_hps_f2h_sdram1_data_awaddr),  //                  .awaddr
		.f2h_sdram1_AWLEN         (mm_interconnect_2_sys_hps_f2h_sdram1_data_awlen),   //                  .awlen
		.f2h_sdram1_AWID          (mm_interconnect_2_sys_hps_f2h_sdram1_data_awid),    //                  .awid
		.f2h_sdram1_AWSIZE        (mm_interconnect_2_sys_hps_f2h_sdram1_data_awsize),  //                  .awsize
		.f2h_sdram1_AWBURST       (mm_interconnect_2_sys_hps_f2h_sdram1_data_awburst), //                  .awburst
		.f2h_sdram1_AWLOCK        (mm_interconnect_2_sys_hps_f2h_sdram1_data_awlock),  //                  .awlock
		.f2h_sdram1_AWPROT        (mm_interconnect_2_sys_hps_f2h_sdram1_data_awprot),  //                  .awprot
		.f2h_sdram1_AWVALID       (mm_interconnect_2_sys_hps_f2h_sdram1_data_awvalid), //                  .awvalid
		.f2h_sdram1_AWCACHE       (mm_interconnect_2_sys_hps_f2h_sdram1_data_awcache), //                  .awcache
		.f2h_sdram1_BRESP         (mm_interconnect_2_sys_hps_f2h_sdram1_data_bresp),   //                  .bresp
		.f2h_sdram1_BID           (mm_interconnect_2_sys_hps_f2h_sdram1_data_bid),     //                  .bid
		.f2h_sdram1_BVALID        (mm_interconnect_2_sys_hps_f2h_sdram1_data_bvalid),  //                  .bvalid
		.f2h_sdram1_BREADY        (mm_interconnect_2_sys_hps_f2h_sdram1_data_bready),  //                  .bready
		.f2h_sdram1_ARREADY       (mm_interconnect_2_sys_hps_f2h_sdram1_data_arready), //                  .arready
		.f2h_sdram1_AWREADY       (mm_interconnect_2_sys_hps_f2h_sdram1_data_awready), //                  .awready
		.f2h_sdram1_RREADY        (mm_interconnect_2_sys_hps_f2h_sdram1_data_rready),  //                  .rready
		.f2h_sdram1_RDATA         (mm_interconnect_2_sys_hps_f2h_sdram1_data_rdata),   //                  .rdata
		.f2h_sdram1_RRESP         (mm_interconnect_2_sys_hps_f2h_sdram1_data_rresp),   //                  .rresp
		.f2h_sdram1_RLAST         (mm_interconnect_2_sys_hps_f2h_sdram1_data_rlast),   //                  .rlast
		.f2h_sdram1_RID           (mm_interconnect_2_sys_hps_f2h_sdram1_data_rid),     //                  .rid
		.f2h_sdram1_RVALID        (mm_interconnect_2_sys_hps_f2h_sdram1_data_rvalid),  //                  .rvalid
		.f2h_sdram1_WLAST         (mm_interconnect_2_sys_hps_f2h_sdram1_data_wlast),   //                  .wlast
		.f2h_sdram1_WVALID        (mm_interconnect_2_sys_hps_f2h_sdram1_data_wvalid),  //                  .wvalid
		.f2h_sdram1_WDATA         (mm_interconnect_2_sys_hps_f2h_sdram1_data_wdata),   //                  .wdata
		.f2h_sdram1_WSTRB         (mm_interconnect_2_sys_hps_f2h_sdram1_data_wstrb),   //                  .wstrb
		.f2h_sdram1_WREADY        (mm_interconnect_2_sys_hps_f2h_sdram1_data_wready),  //                  .wready
		.f2h_sdram1_WID           (mm_interconnect_2_sys_hps_f2h_sdram1_data_wid),     //                  .wid
		.f2h_sdram2_clk           (sys_hps_h2f_user0_clock_clk),                       //  f2h_sdram2_clock.clk
		.f2h_sdram2_ARADDR        (),                                                  //   f2h_sdram2_data.araddr
		.f2h_sdram2_ARLEN         (),                                                  //                  .arlen
		.f2h_sdram2_ARID          (),                                                  //                  .arid
		.f2h_sdram2_ARSIZE        (),                                                  //                  .arsize
		.f2h_sdram2_ARBURST       (),                                                  //                  .arburst
		.f2h_sdram2_ARLOCK        (),                                                  //                  .arlock
		.f2h_sdram2_ARPROT        (),                                                  //                  .arprot
		.f2h_sdram2_ARVALID       (),                                                  //                  .arvalid
		.f2h_sdram2_ARCACHE       (),                                                  //                  .arcache
		.f2h_sdram2_AWADDR        (),                                                  //                  .awaddr
		.f2h_sdram2_AWLEN         (),                                                  //                  .awlen
		.f2h_sdram2_AWID          (),                                                  //                  .awid
		.f2h_sdram2_AWSIZE        (),                                                  //                  .awsize
		.f2h_sdram2_AWBURST       (),                                                  //                  .awburst
		.f2h_sdram2_AWLOCK        (),                                                  //                  .awlock
		.f2h_sdram2_AWPROT        (),                                                  //                  .awprot
		.f2h_sdram2_AWVALID       (),                                                  //                  .awvalid
		.f2h_sdram2_AWCACHE       (),                                                  //                  .awcache
		.f2h_sdram2_BRESP         (),                                                  //                  .bresp
		.f2h_sdram2_BID           (),                                                  //                  .bid
		.f2h_sdram2_BVALID        (),                                                  //                  .bvalid
		.f2h_sdram2_BREADY        (),                                                  //                  .bready
		.f2h_sdram2_ARREADY       (),                                                  //                  .arready
		.f2h_sdram2_AWREADY       (),                                                  //                  .awready
		.f2h_sdram2_RREADY        (),                                                  //                  .rready
		.f2h_sdram2_RDATA         (),                                                  //                  .rdata
		.f2h_sdram2_RRESP         (),                                                  //                  .rresp
		.f2h_sdram2_RLAST         (),                                                  //                  .rlast
		.f2h_sdram2_RID           (),                                                  //                  .rid
		.f2h_sdram2_RVALID        (),                                                  //                  .rvalid
		.f2h_sdram2_WLAST         (),                                                  //                  .wlast
		.f2h_sdram2_WVALID        (),                                                  //                  .wvalid
		.f2h_sdram2_WDATA         (),                                                  //                  .wdata
		.f2h_sdram2_WSTRB         (),                                                  //                  .wstrb
		.f2h_sdram2_WREADY        (),                                                  //                  .wready
		.f2h_sdram2_WID           (),                                                  //                  .wid
		.h2f_axi_clk              (sys_clk_clk),                                       //     h2f_axi_clock.clk
		.h2f_AWID                 (sys_hps_h2f_axi_master_awid),                       //    h2f_axi_master.awid
		.h2f_AWADDR               (sys_hps_h2f_axi_master_awaddr),                     //                  .awaddr
		.h2f_AWLEN                (sys_hps_h2f_axi_master_awlen),                      //                  .awlen
		.h2f_AWSIZE               (sys_hps_h2f_axi_master_awsize),                     //                  .awsize
		.h2f_AWBURST              (sys_hps_h2f_axi_master_awburst),                    //                  .awburst
		.h2f_AWLOCK               (sys_hps_h2f_axi_master_awlock),                     //                  .awlock
		.h2f_AWCACHE              (sys_hps_h2f_axi_master_awcache),                    //                  .awcache
		.h2f_AWPROT               (sys_hps_h2f_axi_master_awprot),                     //                  .awprot
		.h2f_AWVALID              (sys_hps_h2f_axi_master_awvalid),                    //                  .awvalid
		.h2f_AWREADY              (sys_hps_h2f_axi_master_awready),                    //                  .awready
		.h2f_WID                  (sys_hps_h2f_axi_master_wid),                        //                  .wid
		.h2f_WDATA                (sys_hps_h2f_axi_master_wdata),                      //                  .wdata
		.h2f_WSTRB                (sys_hps_h2f_axi_master_wstrb),                      //                  .wstrb
		.h2f_WLAST                (sys_hps_h2f_axi_master_wlast),                      //                  .wlast
		.h2f_WVALID               (sys_hps_h2f_axi_master_wvalid),                     //                  .wvalid
		.h2f_WREADY               (sys_hps_h2f_axi_master_wready),                     //                  .wready
		.h2f_BID                  (sys_hps_h2f_axi_master_bid),                        //                  .bid
		.h2f_BRESP                (sys_hps_h2f_axi_master_bresp),                      //                  .bresp
		.h2f_BVALID               (sys_hps_h2f_axi_master_bvalid),                     //                  .bvalid
		.h2f_BREADY               (sys_hps_h2f_axi_master_bready),                     //                  .bready
		.h2f_ARID                 (sys_hps_h2f_axi_master_arid),                       //                  .arid
		.h2f_ARADDR               (sys_hps_h2f_axi_master_araddr),                     //                  .araddr
		.h2f_ARLEN                (sys_hps_h2f_axi_master_arlen),                      //                  .arlen
		.h2f_ARSIZE               (sys_hps_h2f_axi_master_arsize),                     //                  .arsize
		.h2f_ARBURST              (sys_hps_h2f_axi_master_arburst),                    //                  .arburst
		.h2f_ARLOCK               (sys_hps_h2f_axi_master_arlock),                     //                  .arlock
		.h2f_ARCACHE              (sys_hps_h2f_axi_master_arcache),                    //                  .arcache
		.h2f_ARPROT               (sys_hps_h2f_axi_master_arprot),                     //                  .arprot
		.h2f_ARVALID              (sys_hps_h2f_axi_master_arvalid),                    //                  .arvalid
		.h2f_ARREADY              (sys_hps_h2f_axi_master_arready),                    //                  .arready
		.h2f_RID                  (sys_hps_h2f_axi_master_rid),                        //                  .rid
		.h2f_RDATA                (sys_hps_h2f_axi_master_rdata),                      //                  .rdata
		.h2f_RRESP                (sys_hps_h2f_axi_master_rresp),                      //                  .rresp
		.h2f_RLAST                (sys_hps_h2f_axi_master_rlast),                      //                  .rlast
		.h2f_RVALID               (sys_hps_h2f_axi_master_rvalid),                     //                  .rvalid
		.h2f_RREADY               (sys_hps_h2f_axi_master_rready),                     //                  .rready
		.f2h_axi_clk              (sys_clk_clk),                                       //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                                  //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                                  //                  .awaddr
		.f2h_AWLEN                (),                                                  //                  .awlen
		.f2h_AWSIZE               (),                                                  //                  .awsize
		.f2h_AWBURST              (),                                                  //                  .awburst
		.f2h_AWLOCK               (),                                                  //                  .awlock
		.f2h_AWCACHE              (),                                                  //                  .awcache
		.f2h_AWPROT               (),                                                  //                  .awprot
		.f2h_AWVALID              (),                                                  //                  .awvalid
		.f2h_AWREADY              (),                                                  //                  .awready
		.f2h_AWUSER               (),                                                  //                  .awuser
		.f2h_WID                  (),                                                  //                  .wid
		.f2h_WDATA                (),                                                  //                  .wdata
		.f2h_WSTRB                (),                                                  //                  .wstrb
		.f2h_WLAST                (),                                                  //                  .wlast
		.f2h_WVALID               (),                                                  //                  .wvalid
		.f2h_WREADY               (),                                                  //                  .wready
		.f2h_BID                  (),                                                  //                  .bid
		.f2h_BRESP                (),                                                  //                  .bresp
		.f2h_BVALID               (),                                                  //                  .bvalid
		.f2h_BREADY               (),                                                  //                  .bready
		.f2h_ARID                 (),                                                  //                  .arid
		.f2h_ARADDR               (),                                                  //                  .araddr
		.f2h_ARLEN                (),                                                  //                  .arlen
		.f2h_ARSIZE               (),                                                  //                  .arsize
		.f2h_ARBURST              (),                                                  //                  .arburst
		.f2h_ARLOCK               (),                                                  //                  .arlock
		.f2h_ARCACHE              (),                                                  //                  .arcache
		.f2h_ARPROT               (),                                                  //                  .arprot
		.f2h_ARVALID              (),                                                  //                  .arvalid
		.f2h_ARREADY              (),                                                  //                  .arready
		.f2h_ARUSER               (),                                                  //                  .aruser
		.f2h_RID                  (),                                                  //                  .rid
		.f2h_RDATA                (),                                                  //                  .rdata
		.f2h_RRESP                (),                                                  //                  .rresp
		.f2h_RLAST                (),                                                  //                  .rlast
		.f2h_RVALID               (),                                                  //                  .rvalid
		.f2h_RREADY               (),                                                  //                  .rready
		.h2f_lw_axi_clk           (sys_clk_clk),                                       //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (sys_hps_h2f_lw_axi_master_awid),                    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (sys_hps_h2f_lw_axi_master_awaddr),                  //                  .awaddr
		.h2f_lw_AWLEN             (sys_hps_h2f_lw_axi_master_awlen),                   //                  .awlen
		.h2f_lw_AWSIZE            (sys_hps_h2f_lw_axi_master_awsize),                  //                  .awsize
		.h2f_lw_AWBURST           (sys_hps_h2f_lw_axi_master_awburst),                 //                  .awburst
		.h2f_lw_AWLOCK            (sys_hps_h2f_lw_axi_master_awlock),                  //                  .awlock
		.h2f_lw_AWCACHE           (sys_hps_h2f_lw_axi_master_awcache),                 //                  .awcache
		.h2f_lw_AWPROT            (sys_hps_h2f_lw_axi_master_awprot),                  //                  .awprot
		.h2f_lw_AWVALID           (sys_hps_h2f_lw_axi_master_awvalid),                 //                  .awvalid
		.h2f_lw_AWREADY           (sys_hps_h2f_lw_axi_master_awready),                 //                  .awready
		.h2f_lw_WID               (sys_hps_h2f_lw_axi_master_wid),                     //                  .wid
		.h2f_lw_WDATA             (sys_hps_h2f_lw_axi_master_wdata),                   //                  .wdata
		.h2f_lw_WSTRB             (sys_hps_h2f_lw_axi_master_wstrb),                   //                  .wstrb
		.h2f_lw_WLAST             (sys_hps_h2f_lw_axi_master_wlast),                   //                  .wlast
		.h2f_lw_WVALID            (sys_hps_h2f_lw_axi_master_wvalid),                  //                  .wvalid
		.h2f_lw_WREADY            (sys_hps_h2f_lw_axi_master_wready),                  //                  .wready
		.h2f_lw_BID               (sys_hps_h2f_lw_axi_master_bid),                     //                  .bid
		.h2f_lw_BRESP             (sys_hps_h2f_lw_axi_master_bresp),                   //                  .bresp
		.h2f_lw_BVALID            (sys_hps_h2f_lw_axi_master_bvalid),                  //                  .bvalid
		.h2f_lw_BREADY            (sys_hps_h2f_lw_axi_master_bready),                  //                  .bready
		.h2f_lw_ARID              (sys_hps_h2f_lw_axi_master_arid),                    //                  .arid
		.h2f_lw_ARADDR            (sys_hps_h2f_lw_axi_master_araddr),                  //                  .araddr
		.h2f_lw_ARLEN             (sys_hps_h2f_lw_axi_master_arlen),                   //                  .arlen
		.h2f_lw_ARSIZE            (sys_hps_h2f_lw_axi_master_arsize),                  //                  .arsize
		.h2f_lw_ARBURST           (sys_hps_h2f_lw_axi_master_arburst),                 //                  .arburst
		.h2f_lw_ARLOCK            (sys_hps_h2f_lw_axi_master_arlock),                  //                  .arlock
		.h2f_lw_ARCACHE           (sys_hps_h2f_lw_axi_master_arcache),                 //                  .arcache
		.h2f_lw_ARPROT            (sys_hps_h2f_lw_axi_master_arprot),                  //                  .arprot
		.h2f_lw_ARVALID           (sys_hps_h2f_lw_axi_master_arvalid),                 //                  .arvalid
		.h2f_lw_ARREADY           (sys_hps_h2f_lw_axi_master_arready),                 //                  .arready
		.h2f_lw_RID               (sys_hps_h2f_lw_axi_master_rid),                     //                  .rid
		.h2f_lw_RDATA             (sys_hps_h2f_lw_axi_master_rdata),                   //                  .rdata
		.h2f_lw_RRESP             (sys_hps_h2f_lw_axi_master_rresp),                   //                  .rresp
		.h2f_lw_RLAST             (sys_hps_h2f_lw_axi_master_rlast),                   //                  .rlast
		.h2f_lw_RVALID            (sys_hps_h2f_lw_axi_master_rvalid),                  //                  .rvalid
		.h2f_lw_RREADY            (sys_hps_h2f_lw_axi_master_rready),                  //                  .rready
		.f2h_irq_p0               (sys_hps_f2h_irq0_irq),                              //          f2h_irq0.irq
		.f2h_irq_p1               (sys_hps_f2h_irq1_irq)                               //          f2h_irq1.irq
	);

	system_bd_sys_id sys_id (
		.clock    (sys_clk_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_1_sys_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sys_id_control_slave_address)   //              .address
	);

	system_bd_sys_int_mem sys_int_mem (
		.clk        (sys_clk_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_sys_int_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sys_int_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sys_int_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sys_int_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sys_int_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sys_int_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sys_int_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze     (1'b0)                                         // (terminated)
	);

	system_bd_sys_spi sys_spi (
		.clk           (sys_clk_clk),                                           //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //            reset.reset_n
		.data_from_cpu (mm_interconnect_1_sys_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_1_sys_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_1_sys_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_1_sys_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_1_sys_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_1_sys_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver3_irq),                              //              irq.irq
		.MISO          (sys_spi_MISO),                                          //         external.export
		.MOSI          (sys_spi_MOSI),                                          //                 .export
		.SCLK          (sys_spi_SCLK),                                          //                 .export
		.SS_n          (sys_spi_SS_n)                                           //                 .export
	);

	util_cpack2_impl #(
		.NUM_OF_CHANNELS     (8),
		.SAMPLES_PER_CHANNEL (1),
		.SAMPLE_DATA_WIDTH   (32)
	) util_adc_pack (
		.clk                     (sys_clk_clk),                                                                                                                                                                                                                                                       //                        clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                                                                                                                                                                    //                      reset.reset
		.packed_fifo_wr_en       (util_adc_pack_if_packed_fifo_wr_en_valid),                                                                                                                                                                                                                          //       if_packed_fifo_wr_en.valid
		.packed_fifo_wr_sync     (util_adc_pack_if_packed_fifo_wr_sync_sync),                                                                                                                                                                                                                         //     if_packed_fifo_wr_sync.sync
		.packed_fifo_wr_data     (util_adc_pack_if_packed_fifo_wr_data_data),                                                                                                                                                                                                                         //     if_packed_fifo_wr_data.data
		.packed_fifo_wr_overflow (axi_adc_dma_if_fifo_wr_overflow_ovf),                                                                                                                                                                                                                               // if_packed_fifo_wr_overflow.ovf
		.fifo_wr_overflow        (util_adc_pack_if_fifo_wr_overflow_ovf),                                                                                                                                                                                                                             //        if_fifo_wr_overflow.ovf
		.enable                  ({axi_ltc235x_adc_ch_7_enable,axi_ltc235x_adc_ch_6_enable,axi_ltc235x_adc_ch_5_enable,axi_ltc235x_adc_ch_4_enable,axi_ltc235x_adc_ch_3_enable,axi_ltc235x_adc_ch_2_enable,axi_ltc235x_adc_ch_1_enable,axi_ltc235x_adc_ch_0_enable}),                                 //                   adc_ch_0.enable
		.fifo_wr_en              ({axi_ltc235x_adc_ch_7_valid,axi_ltc235x_adc_ch_6_valid,axi_ltc235x_adc_ch_5_valid,axi_ltc235x_adc_ch_4_valid,axi_ltc235x_adc_ch_3_valid,axi_ltc235x_adc_ch_2_valid,axi_ltc235x_adc_ch_1_valid,axi_ltc235x_adc_ch_0_valid}),                                         //                           .valid
		.fifo_wr_data            ({axi_ltc235x_adc_ch_7_data[31:0],axi_ltc235x_adc_ch_6_data[31:0],axi_ltc235x_adc_ch_5_data[31:0],axi_ltc235x_adc_ch_4_data[31:0],axi_ltc235x_adc_ch_3_data[31:0],axi_ltc235x_adc_ch_2_data[31:0],axi_ltc235x_adc_ch_1_data[31:0],axi_ltc235x_adc_ch_0_data[31:0]})  //                           .data
	);

	axi_hdmi_tx #(
		.ID              (0),
		.CR_CB_N         (0),
		.FPGA_TECHNOLOGY (101)
	) vga_out (
		.s_axi_aclk        (sys_clk_clk),                             //   s_axi_clock.clk
		.s_axi_aresetn     (~rst_controller_reset_out_reset),         //   s_axi_reset.reset_n
		.s_axi_awvalid     (mm_interconnect_1_vga_out_s_axi_awvalid), //         s_axi.awvalid
		.s_axi_awaddr      (mm_interconnect_1_vga_out_s_axi_awaddr),  //              .awaddr
		.s_axi_awprot      (mm_interconnect_1_vga_out_s_axi_awprot),  //              .awprot
		.s_axi_awready     (mm_interconnect_1_vga_out_s_axi_awready), //              .awready
		.s_axi_wvalid      (mm_interconnect_1_vga_out_s_axi_wvalid),  //              .wvalid
		.s_axi_wdata       (mm_interconnect_1_vga_out_s_axi_wdata),   //              .wdata
		.s_axi_wstrb       (mm_interconnect_1_vga_out_s_axi_wstrb),   //              .wstrb
		.s_axi_wready      (mm_interconnect_1_vga_out_s_axi_wready),  //              .wready
		.s_axi_bvalid      (mm_interconnect_1_vga_out_s_axi_bvalid),  //              .bvalid
		.s_axi_bresp       (mm_interconnect_1_vga_out_s_axi_bresp),   //              .bresp
		.s_axi_bready      (mm_interconnect_1_vga_out_s_axi_bready),  //              .bready
		.s_axi_arvalid     (mm_interconnect_1_vga_out_s_axi_arvalid), //              .arvalid
		.s_axi_araddr      (mm_interconnect_1_vga_out_s_axi_araddr),  //              .araddr
		.s_axi_arprot      (mm_interconnect_1_vga_out_s_axi_arprot),  //              .arprot
		.s_axi_arready     (mm_interconnect_1_vga_out_s_axi_arready), //              .arready
		.s_axi_rvalid      (mm_interconnect_1_vga_out_s_axi_rvalid),  //              .rvalid
		.s_axi_rresp       (mm_interconnect_1_vga_out_s_axi_rresp),   //              .rresp
		.s_axi_rdata       (mm_interconnect_1_vga_out_s_axi_rdata),   //              .rdata
		.s_axi_rready      (mm_interconnect_1_vga_out_s_axi_rready),  //              .rready
		.reference_clk     (pixel_clk_pll_outclk0_clk),               // reference_clk.clk
		.vdma_clk          (pixel_clk_pll_outclk1_clk),               //    vdma_clock.clk
		.vdma_valid        (video_dmac_m_axis_tvalid),                //       vdma_if.tvalid
		.vdma_data         (video_dmac_m_axis_tdata),                 //              .tdata
		.vdma_ready        (video_dmac_m_axis_tready),                //              .tready
		.vdma_end_of_frame (video_dmac_m_axis_tlast),                 //              .tlast
		.vga_out_clk       (vga_out_vga_if_vga_clk),                  //        vga_if.vga_clk
		.vga_hsync         (vga_out_vga_if_vga_hsync),                //              .vga_hsync
		.vga_vsync         (vga_out_vga_if_vga_vsync),                //              .vga_vsync
		.vga_red           (vga_out_vga_if_vga_red),                  //              .vga_red
		.vga_green         (vga_out_vga_if_vga_green),                //              .vga_green
		.vga_blue          (vga_out_vga_if_vga_blue)                  //              .vga_blue
	);

	axi_dmac #(
		.ID                    (0),
		.DMA_LENGTH_WIDTH      (24),
		.FIFO_SIZE             (8),
		.MAX_BYTES_PER_BURST   (128),
		.DMA_TYPE_SRC          (0),
		.DMA_AXI_PROTOCOL_SRC  (1),
		.DMA_DATA_WIDTH_SRC    (64),
		.AXI_SLICE_SRC         (0),
		.DMA_TYPE_DEST         (1),
		.DMA_AXI_PROTOCOL_DEST (1),
		.DMA_DATA_WIDTH_DEST   (64),
		.AXI_SLICE_DEST        (0),
		.CYCLIC                (1),
		.DMA_2D_TRANSFER       (1),
		.SYNC_TRANSFER_START   (0),
		.ASYNC_CLK_REQ_SRC     (1),
		.ASYNC_CLK_SRC_DEST    (0),
		.ASYNC_CLK_DEST_REQ    (1),
		.ENABLE_DIAGNOSTICS_IF (0),
		.DMA_AXIS_ID_W         (8),
		.DMA_AXIS_DEST_W       (4)
	) video_dmac (
		.s_axi_aclk             (sys_clk_clk),                                                          //        s_axi_clock.clk
		.s_axi_aresetn          (~rst_controller_reset_out_reset),                                      //        s_axi_reset.reset_n
		.s_axi_awvalid          (mm_interconnect_1_video_dmac_s_axi_awvalid),                           //              s_axi.awvalid
		.s_axi_awaddr           (mm_interconnect_1_video_dmac_s_axi_awaddr),                            //                   .awaddr
		.s_axi_awprot           (mm_interconnect_1_video_dmac_s_axi_awprot),                            //                   .awprot
		.s_axi_awready          (mm_interconnect_1_video_dmac_s_axi_awready),                           //                   .awready
		.s_axi_wvalid           (mm_interconnect_1_video_dmac_s_axi_wvalid),                            //                   .wvalid
		.s_axi_wdata            (mm_interconnect_1_video_dmac_s_axi_wdata),                             //                   .wdata
		.s_axi_wstrb            (mm_interconnect_1_video_dmac_s_axi_wstrb),                             //                   .wstrb
		.s_axi_wready           (mm_interconnect_1_video_dmac_s_axi_wready),                            //                   .wready
		.s_axi_bvalid           (mm_interconnect_1_video_dmac_s_axi_bvalid),                            //                   .bvalid
		.s_axi_bresp            (mm_interconnect_1_video_dmac_s_axi_bresp),                             //                   .bresp
		.s_axi_bready           (mm_interconnect_1_video_dmac_s_axi_bready),                            //                   .bready
		.s_axi_arvalid          (mm_interconnect_1_video_dmac_s_axi_arvalid),                           //                   .arvalid
		.s_axi_araddr           (mm_interconnect_1_video_dmac_s_axi_araddr),                            //                   .araddr
		.s_axi_arprot           (mm_interconnect_1_video_dmac_s_axi_arprot),                            //                   .arprot
		.s_axi_arready          (mm_interconnect_1_video_dmac_s_axi_arready),                           //                   .arready
		.s_axi_rvalid           (mm_interconnect_1_video_dmac_s_axi_rvalid),                            //                   .rvalid
		.s_axi_rresp            (mm_interconnect_1_video_dmac_s_axi_rresp),                             //                   .rresp
		.s_axi_rdata            (mm_interconnect_1_video_dmac_s_axi_rdata),                             //                   .rdata
		.s_axi_rready           (mm_interconnect_1_video_dmac_s_axi_rready),                            //                   .rready
		.irq                    (irq_mapper_receiver0_irq),                                             //   interrupt_sender.irq
		.m_src_axi_aclk         (pixel_clk_pll_outclk1_clk),                                            //    m_src_axi_clock.clk
		.m_src_axi_aresetn      (~rst_controller_001_reset_out_reset),                                  //    m_src_axi_reset.reset_n
		.m_axis_aclk            (pixel_clk_pll_outclk1_clk),                                            //     if_m_axis_aclk.clk
		.m_axis_xfer_req        (),                                                                     // if_m_axis_xfer_req.xfer_req
		.m_axis_valid           (video_dmac_m_axis_tvalid),                                             //             m_axis.tvalid
		.m_axis_last            (video_dmac_m_axis_tlast),                                              //                   .tlast
		.m_axis_ready           (video_dmac_m_axis_tready),                                             //                   .tready
		.m_axis_data            (video_dmac_m_axis_tdata),                                              //                   .tdata
		.m_src_axi_awvalid      (video_dmac_m_src_axi_awvalid),                                         //          m_src_axi.awvalid
		.m_src_axi_awaddr       (video_dmac_m_src_axi_awaddr),                                          //                   .awaddr
		.m_src_axi_awready      (video_dmac_m_src_axi_awready),                                         //                   .awready
		.m_src_axi_wvalid       (video_dmac_m_src_axi_wvalid),                                          //                   .wvalid
		.m_src_axi_wdata        (video_dmac_m_src_axi_wdata),                                           //                   .wdata
		.m_src_axi_wstrb        (video_dmac_m_src_axi_wstrb),                                           //                   .wstrb
		.m_src_axi_wready       (video_dmac_m_src_axi_wready),                                          //                   .wready
		.m_src_axi_bvalid       (video_dmac_m_src_axi_bvalid),                                          //                   .bvalid
		.m_src_axi_bresp        (video_dmac_m_src_axi_bresp),                                           //                   .bresp
		.m_src_axi_bready       (video_dmac_m_src_axi_bready),                                          //                   .bready
		.m_src_axi_arvalid      (video_dmac_m_src_axi_arvalid),                                         //                   .arvalid
		.m_src_axi_araddr       (video_dmac_m_src_axi_araddr),                                          //                   .araddr
		.m_src_axi_arready      (video_dmac_m_src_axi_arready),                                         //                   .arready
		.m_src_axi_rvalid       (video_dmac_m_src_axi_rvalid),                                          //                   .rvalid
		.m_src_axi_rresp        (video_dmac_m_src_axi_rresp),                                           //                   .rresp
		.m_src_axi_rdata        (video_dmac_m_src_axi_rdata),                                           //                   .rdata
		.m_src_axi_rready       (video_dmac_m_src_axi_rready),                                          //                   .rready
		.m_src_axi_awlen        (video_dmac_m_src_axi_awlen),                                           //                   .awlen
		.m_src_axi_awsize       (video_dmac_m_src_axi_awsize),                                          //                   .awsize
		.m_src_axi_awburst      (video_dmac_m_src_axi_awburst),                                         //                   .awburst
		.m_src_axi_awcache      (video_dmac_m_src_axi_awcache),                                         //                   .awcache
		.m_src_axi_awprot       (video_dmac_m_src_axi_awprot),                                          //                   .awprot
		.m_src_axi_wlast        (video_dmac_m_src_axi_wlast),                                           //                   .wlast
		.m_src_axi_arlen        (video_dmac_m_src_axi_arlen),                                           //                   .arlen
		.m_src_axi_arsize       (video_dmac_m_src_axi_arsize),                                          //                   .arsize
		.m_src_axi_arburst      (video_dmac_m_src_axi_arburst),                                         //                   .arburst
		.m_src_axi_arcache      (video_dmac_m_src_axi_arcache),                                         //                   .arcache
		.m_src_axi_arprot       (video_dmac_m_src_axi_arprot),                                          //                   .arprot
		.m_src_axi_awid         (video_dmac_m_src_axi_awid),                                            //                   .awid
		.m_src_axi_awlock       (video_dmac_m_src_axi_awlock),                                          //                   .awlock
		.m_src_axi_wid          (video_dmac_m_src_axi_wid),                                             //                   .wid
		.m_src_axi_arid         (video_dmac_m_src_axi_arid),                                            //                   .arid
		.m_src_axi_arlock       (video_dmac_m_src_axi_arlock),                                          //                   .arlock
		.m_src_axi_rid          (video_dmac_m_src_axi_rid),                                             //                   .rid
		.m_src_axi_bid          (video_dmac_m_src_axi_bid),                                             //                   .bid
		.m_src_axi_rlast        (video_dmac_m_src_axi_rlast),                                           //                   .rlast
		.m_axis_user            (),                                                                     //        (terminated)
		.m_axis_id              (),                                                                     //        (terminated)
		.m_axis_dest            (),                                                                     //        (terminated)
		.m_axis_strb            (),                                                                     //        (terminated)
		.m_axis_keep            (),                                                                     //        (terminated)
		.m_dest_axi_aclk        (1'b0),                                                                 //        (terminated)
		.m_dest_axi_aresetn     (1'b1),                                                                 //        (terminated)
		.s_axis_aclk            (1'b0),                                                                 //        (terminated)
		.s_axis_xfer_req        (),                                                                     //        (terminated)
		.s_axis_valid           (1'b0),                                                                 //        (terminated)
		.s_axis_last            (1'b0),                                                                 //        (terminated)
		.s_axis_ready           (),                                                                     //        (terminated)
		.s_axis_data            (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.s_axis_user            (1'b0),                                                                 //        (terminated)
		.s_axis_id              (8'b00000000),                                                          //        (terminated)
		.s_axis_dest            (4'b0000),                                                              //        (terminated)
		.s_axis_strb            (8'b00000000),                                                          //        (terminated)
		.s_axis_keep            (8'b00000000),                                                          //        (terminated)
		.fifo_rd_clk            (1'b0),                                                                 //        (terminated)
		.fifo_rd_en             (1'b0),                                                                 //        (terminated)
		.fifo_rd_valid          (),                                                                     //        (terminated)
		.fifo_rd_dout           (),                                                                     //        (terminated)
		.fifo_rd_underflow      (),                                                                     //        (terminated)
		.fifo_rd_xfer_req       (),                                                                     //        (terminated)
		.fifo_wr_clk            (1'b0),                                                                 //        (terminated)
		.fifo_wr_en             (1'b0),                                                                 //        (terminated)
		.fifo_wr_din            (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.fifo_wr_overflow       (),                                                                     //        (terminated)
		.fifo_wr_sync           (1'b0),                                                                 //        (terminated)
		.fifo_wr_xfer_req       (),                                                                     //        (terminated)
		.dest_diag_level_bursts (),                                                                     //        (terminated)
		.m_dest_axi_awvalid     (),                                                                     //        (terminated)
		.m_dest_axi_awaddr      (),                                                                     //        (terminated)
		.m_dest_axi_awready     (1'b0),                                                                 //        (terminated)
		.m_dest_axi_wvalid      (),                                                                     //        (terminated)
		.m_dest_axi_wdata       (),                                                                     //        (terminated)
		.m_dest_axi_wstrb       (),                                                                     //        (terminated)
		.m_dest_axi_wready      (1'b0),                                                                 //        (terminated)
		.m_dest_axi_bvalid      (1'b0),                                                                 //        (terminated)
		.m_dest_axi_bresp       (2'b00),                                                                //        (terminated)
		.m_dest_axi_bready      (),                                                                     //        (terminated)
		.m_dest_axi_arvalid     (),                                                                     //        (terminated)
		.m_dest_axi_araddr      (),                                                                     //        (terminated)
		.m_dest_axi_arready     (1'b0),                                                                 //        (terminated)
		.m_dest_axi_rvalid      (1'b0),                                                                 //        (terminated)
		.m_dest_axi_rresp       (2'b00),                                                                //        (terminated)
		.m_dest_axi_rdata       (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.m_dest_axi_rready      (),                                                                     //        (terminated)
		.m_dest_axi_awlen       (),                                                                     //        (terminated)
		.m_dest_axi_awsize      (),                                                                     //        (terminated)
		.m_dest_axi_awburst     (),                                                                     //        (terminated)
		.m_dest_axi_awcache     (),                                                                     //        (terminated)
		.m_dest_axi_awprot      (),                                                                     //        (terminated)
		.m_dest_axi_wlast       (),                                                                     //        (terminated)
		.m_dest_axi_arlen       (),                                                                     //        (terminated)
		.m_dest_axi_arsize      (),                                                                     //        (terminated)
		.m_dest_axi_arburst     (),                                                                     //        (terminated)
		.m_dest_axi_arcache     (),                                                                     //        (terminated)
		.m_dest_axi_arprot      (),                                                                     //        (terminated)
		.m_dest_axi_awid        (),                                                                     //        (terminated)
		.m_dest_axi_awlock      (),                                                                     //        (terminated)
		.m_dest_axi_wid         (),                                                                     //        (terminated)
		.m_dest_axi_arid        (),                                                                     //        (terminated)
		.m_dest_axi_arlock      (),                                                                     //        (terminated)
		.m_dest_axi_rid         (1'b0),                                                                 //        (terminated)
		.m_dest_axi_bid         (1'b0),                                                                 //        (terminated)
		.m_dest_axi_rlast       (1'b0)                                                                  //        (terminated)
	);

	system_bd_mm_interconnect_0 mm_interconnect_0 (
		.sys_hps_h2f_axi_master_awid                                        (sys_hps_h2f_axi_master_awid),                 //                                       sys_hps_h2f_axi_master.awid
		.sys_hps_h2f_axi_master_awaddr                                      (sys_hps_h2f_axi_master_awaddr),               //                                                             .awaddr
		.sys_hps_h2f_axi_master_awlen                                       (sys_hps_h2f_axi_master_awlen),                //                                                             .awlen
		.sys_hps_h2f_axi_master_awsize                                      (sys_hps_h2f_axi_master_awsize),               //                                                             .awsize
		.sys_hps_h2f_axi_master_awburst                                     (sys_hps_h2f_axi_master_awburst),              //                                                             .awburst
		.sys_hps_h2f_axi_master_awlock                                      (sys_hps_h2f_axi_master_awlock),               //                                                             .awlock
		.sys_hps_h2f_axi_master_awcache                                     (sys_hps_h2f_axi_master_awcache),              //                                                             .awcache
		.sys_hps_h2f_axi_master_awprot                                      (sys_hps_h2f_axi_master_awprot),               //                                                             .awprot
		.sys_hps_h2f_axi_master_awvalid                                     (sys_hps_h2f_axi_master_awvalid),              //                                                             .awvalid
		.sys_hps_h2f_axi_master_awready                                     (sys_hps_h2f_axi_master_awready),              //                                                             .awready
		.sys_hps_h2f_axi_master_wid                                         (sys_hps_h2f_axi_master_wid),                  //                                                             .wid
		.sys_hps_h2f_axi_master_wdata                                       (sys_hps_h2f_axi_master_wdata),                //                                                             .wdata
		.sys_hps_h2f_axi_master_wstrb                                       (sys_hps_h2f_axi_master_wstrb),                //                                                             .wstrb
		.sys_hps_h2f_axi_master_wlast                                       (sys_hps_h2f_axi_master_wlast),                //                                                             .wlast
		.sys_hps_h2f_axi_master_wvalid                                      (sys_hps_h2f_axi_master_wvalid),               //                                                             .wvalid
		.sys_hps_h2f_axi_master_wready                                      (sys_hps_h2f_axi_master_wready),               //                                                             .wready
		.sys_hps_h2f_axi_master_bid                                         (sys_hps_h2f_axi_master_bid),                  //                                                             .bid
		.sys_hps_h2f_axi_master_bresp                                       (sys_hps_h2f_axi_master_bresp),                //                                                             .bresp
		.sys_hps_h2f_axi_master_bvalid                                      (sys_hps_h2f_axi_master_bvalid),               //                                                             .bvalid
		.sys_hps_h2f_axi_master_bready                                      (sys_hps_h2f_axi_master_bready),               //                                                             .bready
		.sys_hps_h2f_axi_master_arid                                        (sys_hps_h2f_axi_master_arid),                 //                                                             .arid
		.sys_hps_h2f_axi_master_araddr                                      (sys_hps_h2f_axi_master_araddr),               //                                                             .araddr
		.sys_hps_h2f_axi_master_arlen                                       (sys_hps_h2f_axi_master_arlen),                //                                                             .arlen
		.sys_hps_h2f_axi_master_arsize                                      (sys_hps_h2f_axi_master_arsize),               //                                                             .arsize
		.sys_hps_h2f_axi_master_arburst                                     (sys_hps_h2f_axi_master_arburst),              //                                                             .arburst
		.sys_hps_h2f_axi_master_arlock                                      (sys_hps_h2f_axi_master_arlock),               //                                                             .arlock
		.sys_hps_h2f_axi_master_arcache                                     (sys_hps_h2f_axi_master_arcache),              //                                                             .arcache
		.sys_hps_h2f_axi_master_arprot                                      (sys_hps_h2f_axi_master_arprot),               //                                                             .arprot
		.sys_hps_h2f_axi_master_arvalid                                     (sys_hps_h2f_axi_master_arvalid),              //                                                             .arvalid
		.sys_hps_h2f_axi_master_arready                                     (sys_hps_h2f_axi_master_arready),              //                                                             .arready
		.sys_hps_h2f_axi_master_rid                                         (sys_hps_h2f_axi_master_rid),                  //                                                             .rid
		.sys_hps_h2f_axi_master_rdata                                       (sys_hps_h2f_axi_master_rdata),                //                                                             .rdata
		.sys_hps_h2f_axi_master_rresp                                       (sys_hps_h2f_axi_master_rresp),                //                                                             .rresp
		.sys_hps_h2f_axi_master_rlast                                       (sys_hps_h2f_axi_master_rlast),                //                                                             .rlast
		.sys_hps_h2f_axi_master_rvalid                                      (sys_hps_h2f_axi_master_rvalid),               //                                                             .rvalid
		.sys_hps_h2f_axi_master_rready                                      (sys_hps_h2f_axi_master_rready),               //                                                             .rready
		.sys_clk_clk_clk                                                    (sys_clk_clk),                                 //                                                  sys_clk_clk.clk
		.sys_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),          // sys_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.sys_int_mem_reset1_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),              //                     sys_int_mem_reset1_reset_bridge_in_reset.reset
		.sys_int_mem_s1_address                                             (mm_interconnect_0_sys_int_mem_s1_address),    //                                               sys_int_mem_s1.address
		.sys_int_mem_s1_write                                               (mm_interconnect_0_sys_int_mem_s1_write),      //                                                             .write
		.sys_int_mem_s1_readdata                                            (mm_interconnect_0_sys_int_mem_s1_readdata),   //                                                             .readdata
		.sys_int_mem_s1_writedata                                           (mm_interconnect_0_sys_int_mem_s1_writedata),  //                                                             .writedata
		.sys_int_mem_s1_byteenable                                          (mm_interconnect_0_sys_int_mem_s1_byteenable), //                                                             .byteenable
		.sys_int_mem_s1_chipselect                                          (mm_interconnect_0_sys_int_mem_s1_chipselect), //                                                             .chipselect
		.sys_int_mem_s1_clken                                               (mm_interconnect_0_sys_int_mem_s1_clken)       //                                                             .clken
	);

	system_bd_mm_interconnect_1 mm_interconnect_1 (
		.adc_pwm_gen_s_axi_awaddr                                              (mm_interconnect_1_adc_pwm_gen_s_axi_awaddr),                             //                                               adc_pwm_gen_s_axi.awaddr
		.adc_pwm_gen_s_axi_awprot                                              (mm_interconnect_1_adc_pwm_gen_s_axi_awprot),                             //                                                                .awprot
		.adc_pwm_gen_s_axi_awvalid                                             (mm_interconnect_1_adc_pwm_gen_s_axi_awvalid),                            //                                                                .awvalid
		.adc_pwm_gen_s_axi_awready                                             (mm_interconnect_1_adc_pwm_gen_s_axi_awready),                            //                                                                .awready
		.adc_pwm_gen_s_axi_wdata                                               (mm_interconnect_1_adc_pwm_gen_s_axi_wdata),                              //                                                                .wdata
		.adc_pwm_gen_s_axi_wstrb                                               (mm_interconnect_1_adc_pwm_gen_s_axi_wstrb),                              //                                                                .wstrb
		.adc_pwm_gen_s_axi_wvalid                                              (mm_interconnect_1_adc_pwm_gen_s_axi_wvalid),                             //                                                                .wvalid
		.adc_pwm_gen_s_axi_wready                                              (mm_interconnect_1_adc_pwm_gen_s_axi_wready),                             //                                                                .wready
		.adc_pwm_gen_s_axi_bresp                                               (mm_interconnect_1_adc_pwm_gen_s_axi_bresp),                              //                                                                .bresp
		.adc_pwm_gen_s_axi_bvalid                                              (mm_interconnect_1_adc_pwm_gen_s_axi_bvalid),                             //                                                                .bvalid
		.adc_pwm_gen_s_axi_bready                                              (mm_interconnect_1_adc_pwm_gen_s_axi_bready),                             //                                                                .bready
		.adc_pwm_gen_s_axi_araddr                                              (mm_interconnect_1_adc_pwm_gen_s_axi_araddr),                             //                                                                .araddr
		.adc_pwm_gen_s_axi_arprot                                              (mm_interconnect_1_adc_pwm_gen_s_axi_arprot),                             //                                                                .arprot
		.adc_pwm_gen_s_axi_arvalid                                             (mm_interconnect_1_adc_pwm_gen_s_axi_arvalid),                            //                                                                .arvalid
		.adc_pwm_gen_s_axi_arready                                             (mm_interconnect_1_adc_pwm_gen_s_axi_arready),                            //                                                                .arready
		.adc_pwm_gen_s_axi_rdata                                               (mm_interconnect_1_adc_pwm_gen_s_axi_rdata),                              //                                                                .rdata
		.adc_pwm_gen_s_axi_rresp                                               (mm_interconnect_1_adc_pwm_gen_s_axi_rresp),                              //                                                                .rresp
		.adc_pwm_gen_s_axi_rvalid                                              (mm_interconnect_1_adc_pwm_gen_s_axi_rvalid),                             //                                                                .rvalid
		.adc_pwm_gen_s_axi_rready                                              (mm_interconnect_1_adc_pwm_gen_s_axi_rready),                             //                                                                .rready
		.axi_adc_dma_s_axi_awaddr                                              (mm_interconnect_1_axi_adc_dma_s_axi_awaddr),                             //                                               axi_adc_dma_s_axi.awaddr
		.axi_adc_dma_s_axi_awprot                                              (mm_interconnect_1_axi_adc_dma_s_axi_awprot),                             //                                                                .awprot
		.axi_adc_dma_s_axi_awvalid                                             (mm_interconnect_1_axi_adc_dma_s_axi_awvalid),                            //                                                                .awvalid
		.axi_adc_dma_s_axi_awready                                             (mm_interconnect_1_axi_adc_dma_s_axi_awready),                            //                                                                .awready
		.axi_adc_dma_s_axi_wdata                                               (mm_interconnect_1_axi_adc_dma_s_axi_wdata),                              //                                                                .wdata
		.axi_adc_dma_s_axi_wstrb                                               (mm_interconnect_1_axi_adc_dma_s_axi_wstrb),                              //                                                                .wstrb
		.axi_adc_dma_s_axi_wvalid                                              (mm_interconnect_1_axi_adc_dma_s_axi_wvalid),                             //                                                                .wvalid
		.axi_adc_dma_s_axi_wready                                              (mm_interconnect_1_axi_adc_dma_s_axi_wready),                             //                                                                .wready
		.axi_adc_dma_s_axi_bresp                                               (mm_interconnect_1_axi_adc_dma_s_axi_bresp),                              //                                                                .bresp
		.axi_adc_dma_s_axi_bvalid                                              (mm_interconnect_1_axi_adc_dma_s_axi_bvalid),                             //                                                                .bvalid
		.axi_adc_dma_s_axi_bready                                              (mm_interconnect_1_axi_adc_dma_s_axi_bready),                             //                                                                .bready
		.axi_adc_dma_s_axi_araddr                                              (mm_interconnect_1_axi_adc_dma_s_axi_araddr),                             //                                                                .araddr
		.axi_adc_dma_s_axi_arprot                                              (mm_interconnect_1_axi_adc_dma_s_axi_arprot),                             //                                                                .arprot
		.axi_adc_dma_s_axi_arvalid                                             (mm_interconnect_1_axi_adc_dma_s_axi_arvalid),                            //                                                                .arvalid
		.axi_adc_dma_s_axi_arready                                             (mm_interconnect_1_axi_adc_dma_s_axi_arready),                            //                                                                .arready
		.axi_adc_dma_s_axi_rdata                                               (mm_interconnect_1_axi_adc_dma_s_axi_rdata),                              //                                                                .rdata
		.axi_adc_dma_s_axi_rresp                                               (mm_interconnect_1_axi_adc_dma_s_axi_rresp),                              //                                                                .rresp
		.axi_adc_dma_s_axi_rvalid                                              (mm_interconnect_1_axi_adc_dma_s_axi_rvalid),                             //                                                                .rvalid
		.axi_adc_dma_s_axi_rready                                              (mm_interconnect_1_axi_adc_dma_s_axi_rready),                             //                                                                .rready
		.axi_ltc235x_s_axi_awaddr                                              (mm_interconnect_1_axi_ltc235x_s_axi_awaddr),                             //                                               axi_ltc235x_s_axi.awaddr
		.axi_ltc235x_s_axi_awprot                                              (mm_interconnect_1_axi_ltc235x_s_axi_awprot),                             //                                                                .awprot
		.axi_ltc235x_s_axi_awvalid                                             (mm_interconnect_1_axi_ltc235x_s_axi_awvalid),                            //                                                                .awvalid
		.axi_ltc235x_s_axi_awready                                             (mm_interconnect_1_axi_ltc235x_s_axi_awready),                            //                                                                .awready
		.axi_ltc235x_s_axi_wdata                                               (mm_interconnect_1_axi_ltc235x_s_axi_wdata),                              //                                                                .wdata
		.axi_ltc235x_s_axi_wstrb                                               (mm_interconnect_1_axi_ltc235x_s_axi_wstrb),                              //                                                                .wstrb
		.axi_ltc235x_s_axi_wvalid                                              (mm_interconnect_1_axi_ltc235x_s_axi_wvalid),                             //                                                                .wvalid
		.axi_ltc235x_s_axi_wready                                              (mm_interconnect_1_axi_ltc235x_s_axi_wready),                             //                                                                .wready
		.axi_ltc235x_s_axi_bresp                                               (mm_interconnect_1_axi_ltc235x_s_axi_bresp),                              //                                                                .bresp
		.axi_ltc235x_s_axi_bvalid                                              (mm_interconnect_1_axi_ltc235x_s_axi_bvalid),                             //                                                                .bvalid
		.axi_ltc235x_s_axi_bready                                              (mm_interconnect_1_axi_ltc235x_s_axi_bready),                             //                                                                .bready
		.axi_ltc235x_s_axi_araddr                                              (mm_interconnect_1_axi_ltc235x_s_axi_araddr),                             //                                                                .araddr
		.axi_ltc235x_s_axi_arprot                                              (mm_interconnect_1_axi_ltc235x_s_axi_arprot),                             //                                                                .arprot
		.axi_ltc235x_s_axi_arvalid                                             (mm_interconnect_1_axi_ltc235x_s_axi_arvalid),                            //                                                                .arvalid
		.axi_ltc235x_s_axi_arready                                             (mm_interconnect_1_axi_ltc235x_s_axi_arready),                            //                                                                .arready
		.axi_ltc235x_s_axi_rdata                                               (mm_interconnect_1_axi_ltc235x_s_axi_rdata),                              //                                                                .rdata
		.axi_ltc235x_s_axi_rresp                                               (mm_interconnect_1_axi_ltc235x_s_axi_rresp),                              //                                                                .rresp
		.axi_ltc235x_s_axi_rvalid                                              (mm_interconnect_1_axi_ltc235x_s_axi_rvalid),                             //                                                                .rvalid
		.axi_ltc235x_s_axi_rready                                              (mm_interconnect_1_axi_ltc235x_s_axi_rready),                             //                                                                .rready
		.axi_sysid_0_s_axi_awaddr                                              (mm_interconnect_1_axi_sysid_0_s_axi_awaddr),                             //                                               axi_sysid_0_s_axi.awaddr
		.axi_sysid_0_s_axi_awprot                                              (mm_interconnect_1_axi_sysid_0_s_axi_awprot),                             //                                                                .awprot
		.axi_sysid_0_s_axi_awvalid                                             (mm_interconnect_1_axi_sysid_0_s_axi_awvalid),                            //                                                                .awvalid
		.axi_sysid_0_s_axi_awready                                             (mm_interconnect_1_axi_sysid_0_s_axi_awready),                            //                                                                .awready
		.axi_sysid_0_s_axi_wdata                                               (mm_interconnect_1_axi_sysid_0_s_axi_wdata),                              //                                                                .wdata
		.axi_sysid_0_s_axi_wstrb                                               (mm_interconnect_1_axi_sysid_0_s_axi_wstrb),                              //                                                                .wstrb
		.axi_sysid_0_s_axi_wvalid                                              (mm_interconnect_1_axi_sysid_0_s_axi_wvalid),                             //                                                                .wvalid
		.axi_sysid_0_s_axi_wready                                              (mm_interconnect_1_axi_sysid_0_s_axi_wready),                             //                                                                .wready
		.axi_sysid_0_s_axi_bresp                                               (mm_interconnect_1_axi_sysid_0_s_axi_bresp),                              //                                                                .bresp
		.axi_sysid_0_s_axi_bvalid                                              (mm_interconnect_1_axi_sysid_0_s_axi_bvalid),                             //                                                                .bvalid
		.axi_sysid_0_s_axi_bready                                              (mm_interconnect_1_axi_sysid_0_s_axi_bready),                             //                                                                .bready
		.axi_sysid_0_s_axi_araddr                                              (mm_interconnect_1_axi_sysid_0_s_axi_araddr),                             //                                                                .araddr
		.axi_sysid_0_s_axi_arprot                                              (mm_interconnect_1_axi_sysid_0_s_axi_arprot),                             //                                                                .arprot
		.axi_sysid_0_s_axi_arvalid                                             (mm_interconnect_1_axi_sysid_0_s_axi_arvalid),                            //                                                                .arvalid
		.axi_sysid_0_s_axi_arready                                             (mm_interconnect_1_axi_sysid_0_s_axi_arready),                            //                                                                .arready
		.axi_sysid_0_s_axi_rdata                                               (mm_interconnect_1_axi_sysid_0_s_axi_rdata),                              //                                                                .rdata
		.axi_sysid_0_s_axi_rresp                                               (mm_interconnect_1_axi_sysid_0_s_axi_rresp),                              //                                                                .rresp
		.axi_sysid_0_s_axi_rvalid                                              (mm_interconnect_1_axi_sysid_0_s_axi_rvalid),                             //                                                                .rvalid
		.axi_sysid_0_s_axi_rready                                              (mm_interconnect_1_axi_sysid_0_s_axi_rready),                             //                                                                .rready
		.sys_hps_h2f_lw_axi_master_awid                                        (sys_hps_h2f_lw_axi_master_awid),                                         //                                       sys_hps_h2f_lw_axi_master.awid
		.sys_hps_h2f_lw_axi_master_awaddr                                      (sys_hps_h2f_lw_axi_master_awaddr),                                       //                                                                .awaddr
		.sys_hps_h2f_lw_axi_master_awlen                                       (sys_hps_h2f_lw_axi_master_awlen),                                        //                                                                .awlen
		.sys_hps_h2f_lw_axi_master_awsize                                      (sys_hps_h2f_lw_axi_master_awsize),                                       //                                                                .awsize
		.sys_hps_h2f_lw_axi_master_awburst                                     (sys_hps_h2f_lw_axi_master_awburst),                                      //                                                                .awburst
		.sys_hps_h2f_lw_axi_master_awlock                                      (sys_hps_h2f_lw_axi_master_awlock),                                       //                                                                .awlock
		.sys_hps_h2f_lw_axi_master_awcache                                     (sys_hps_h2f_lw_axi_master_awcache),                                      //                                                                .awcache
		.sys_hps_h2f_lw_axi_master_awprot                                      (sys_hps_h2f_lw_axi_master_awprot),                                       //                                                                .awprot
		.sys_hps_h2f_lw_axi_master_awvalid                                     (sys_hps_h2f_lw_axi_master_awvalid),                                      //                                                                .awvalid
		.sys_hps_h2f_lw_axi_master_awready                                     (sys_hps_h2f_lw_axi_master_awready),                                      //                                                                .awready
		.sys_hps_h2f_lw_axi_master_wid                                         (sys_hps_h2f_lw_axi_master_wid),                                          //                                                                .wid
		.sys_hps_h2f_lw_axi_master_wdata                                       (sys_hps_h2f_lw_axi_master_wdata),                                        //                                                                .wdata
		.sys_hps_h2f_lw_axi_master_wstrb                                       (sys_hps_h2f_lw_axi_master_wstrb),                                        //                                                                .wstrb
		.sys_hps_h2f_lw_axi_master_wlast                                       (sys_hps_h2f_lw_axi_master_wlast),                                        //                                                                .wlast
		.sys_hps_h2f_lw_axi_master_wvalid                                      (sys_hps_h2f_lw_axi_master_wvalid),                                       //                                                                .wvalid
		.sys_hps_h2f_lw_axi_master_wready                                      (sys_hps_h2f_lw_axi_master_wready),                                       //                                                                .wready
		.sys_hps_h2f_lw_axi_master_bid                                         (sys_hps_h2f_lw_axi_master_bid),                                          //                                                                .bid
		.sys_hps_h2f_lw_axi_master_bresp                                       (sys_hps_h2f_lw_axi_master_bresp),                                        //                                                                .bresp
		.sys_hps_h2f_lw_axi_master_bvalid                                      (sys_hps_h2f_lw_axi_master_bvalid),                                       //                                                                .bvalid
		.sys_hps_h2f_lw_axi_master_bready                                      (sys_hps_h2f_lw_axi_master_bready),                                       //                                                                .bready
		.sys_hps_h2f_lw_axi_master_arid                                        (sys_hps_h2f_lw_axi_master_arid),                                         //                                                                .arid
		.sys_hps_h2f_lw_axi_master_araddr                                      (sys_hps_h2f_lw_axi_master_araddr),                                       //                                                                .araddr
		.sys_hps_h2f_lw_axi_master_arlen                                       (sys_hps_h2f_lw_axi_master_arlen),                                        //                                                                .arlen
		.sys_hps_h2f_lw_axi_master_arsize                                      (sys_hps_h2f_lw_axi_master_arsize),                                       //                                                                .arsize
		.sys_hps_h2f_lw_axi_master_arburst                                     (sys_hps_h2f_lw_axi_master_arburst),                                      //                                                                .arburst
		.sys_hps_h2f_lw_axi_master_arlock                                      (sys_hps_h2f_lw_axi_master_arlock),                                       //                                                                .arlock
		.sys_hps_h2f_lw_axi_master_arcache                                     (sys_hps_h2f_lw_axi_master_arcache),                                      //                                                                .arcache
		.sys_hps_h2f_lw_axi_master_arprot                                      (sys_hps_h2f_lw_axi_master_arprot),                                       //                                                                .arprot
		.sys_hps_h2f_lw_axi_master_arvalid                                     (sys_hps_h2f_lw_axi_master_arvalid),                                      //                                                                .arvalid
		.sys_hps_h2f_lw_axi_master_arready                                     (sys_hps_h2f_lw_axi_master_arready),                                      //                                                                .arready
		.sys_hps_h2f_lw_axi_master_rid                                         (sys_hps_h2f_lw_axi_master_rid),                                          //                                                                .rid
		.sys_hps_h2f_lw_axi_master_rdata                                       (sys_hps_h2f_lw_axi_master_rdata),                                        //                                                                .rdata
		.sys_hps_h2f_lw_axi_master_rresp                                       (sys_hps_h2f_lw_axi_master_rresp),                                        //                                                                .rresp
		.sys_hps_h2f_lw_axi_master_rlast                                       (sys_hps_h2f_lw_axi_master_rlast),                                        //                                                                .rlast
		.sys_hps_h2f_lw_axi_master_rvalid                                      (sys_hps_h2f_lw_axi_master_rvalid),                                       //                                                                .rvalid
		.sys_hps_h2f_lw_axi_master_rready                                      (sys_hps_h2f_lw_axi_master_rready),                                       //                                                                .rready
		.vga_out_s_axi_awaddr                                                  (mm_interconnect_1_vga_out_s_axi_awaddr),                                 //                                                   vga_out_s_axi.awaddr
		.vga_out_s_axi_awprot                                                  (mm_interconnect_1_vga_out_s_axi_awprot),                                 //                                                                .awprot
		.vga_out_s_axi_awvalid                                                 (mm_interconnect_1_vga_out_s_axi_awvalid),                                //                                                                .awvalid
		.vga_out_s_axi_awready                                                 (mm_interconnect_1_vga_out_s_axi_awready),                                //                                                                .awready
		.vga_out_s_axi_wdata                                                   (mm_interconnect_1_vga_out_s_axi_wdata),                                  //                                                                .wdata
		.vga_out_s_axi_wstrb                                                   (mm_interconnect_1_vga_out_s_axi_wstrb),                                  //                                                                .wstrb
		.vga_out_s_axi_wvalid                                                  (mm_interconnect_1_vga_out_s_axi_wvalid),                                 //                                                                .wvalid
		.vga_out_s_axi_wready                                                  (mm_interconnect_1_vga_out_s_axi_wready),                                 //                                                                .wready
		.vga_out_s_axi_bresp                                                   (mm_interconnect_1_vga_out_s_axi_bresp),                                  //                                                                .bresp
		.vga_out_s_axi_bvalid                                                  (mm_interconnect_1_vga_out_s_axi_bvalid),                                 //                                                                .bvalid
		.vga_out_s_axi_bready                                                  (mm_interconnect_1_vga_out_s_axi_bready),                                 //                                                                .bready
		.vga_out_s_axi_araddr                                                  (mm_interconnect_1_vga_out_s_axi_araddr),                                 //                                                                .araddr
		.vga_out_s_axi_arprot                                                  (mm_interconnect_1_vga_out_s_axi_arprot),                                 //                                                                .arprot
		.vga_out_s_axi_arvalid                                                 (mm_interconnect_1_vga_out_s_axi_arvalid),                                //                                                                .arvalid
		.vga_out_s_axi_arready                                                 (mm_interconnect_1_vga_out_s_axi_arready),                                //                                                                .arready
		.vga_out_s_axi_rdata                                                   (mm_interconnect_1_vga_out_s_axi_rdata),                                  //                                                                .rdata
		.vga_out_s_axi_rresp                                                   (mm_interconnect_1_vga_out_s_axi_rresp),                                  //                                                                .rresp
		.vga_out_s_axi_rvalid                                                  (mm_interconnect_1_vga_out_s_axi_rvalid),                                 //                                                                .rvalid
		.vga_out_s_axi_rready                                                  (mm_interconnect_1_vga_out_s_axi_rready),                                 //                                                                .rready
		.video_dmac_s_axi_awaddr                                               (mm_interconnect_1_video_dmac_s_axi_awaddr),                              //                                                video_dmac_s_axi.awaddr
		.video_dmac_s_axi_awprot                                               (mm_interconnect_1_video_dmac_s_axi_awprot),                              //                                                                .awprot
		.video_dmac_s_axi_awvalid                                              (mm_interconnect_1_video_dmac_s_axi_awvalid),                             //                                                                .awvalid
		.video_dmac_s_axi_awready                                              (mm_interconnect_1_video_dmac_s_axi_awready),                             //                                                                .awready
		.video_dmac_s_axi_wdata                                                (mm_interconnect_1_video_dmac_s_axi_wdata),                               //                                                                .wdata
		.video_dmac_s_axi_wstrb                                                (mm_interconnect_1_video_dmac_s_axi_wstrb),                               //                                                                .wstrb
		.video_dmac_s_axi_wvalid                                               (mm_interconnect_1_video_dmac_s_axi_wvalid),                              //                                                                .wvalid
		.video_dmac_s_axi_wready                                               (mm_interconnect_1_video_dmac_s_axi_wready),                              //                                                                .wready
		.video_dmac_s_axi_bresp                                                (mm_interconnect_1_video_dmac_s_axi_bresp),                               //                                                                .bresp
		.video_dmac_s_axi_bvalid                                               (mm_interconnect_1_video_dmac_s_axi_bvalid),                              //                                                                .bvalid
		.video_dmac_s_axi_bready                                               (mm_interconnect_1_video_dmac_s_axi_bready),                              //                                                                .bready
		.video_dmac_s_axi_araddr                                               (mm_interconnect_1_video_dmac_s_axi_araddr),                              //                                                                .araddr
		.video_dmac_s_axi_arprot                                               (mm_interconnect_1_video_dmac_s_axi_arprot),                              //                                                                .arprot
		.video_dmac_s_axi_arvalid                                              (mm_interconnect_1_video_dmac_s_axi_arvalid),                             //                                                                .arvalid
		.video_dmac_s_axi_arready                                              (mm_interconnect_1_video_dmac_s_axi_arready),                             //                                                                .arready
		.video_dmac_s_axi_rdata                                                (mm_interconnect_1_video_dmac_s_axi_rdata),                               //                                                                .rdata
		.video_dmac_s_axi_rresp                                                (mm_interconnect_1_video_dmac_s_axi_rresp),                               //                                                                .rresp
		.video_dmac_s_axi_rvalid                                               (mm_interconnect_1_video_dmac_s_axi_rvalid),                              //                                                                .rvalid
		.video_dmac_s_axi_rready                                               (mm_interconnect_1_video_dmac_s_axi_rready),                              //                                                                .rready
		.sys_clk_clk_clk                                                       (sys_clk_clk),                                                            //                                                     sys_clk_clk.clk
		.sys_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                     // sys_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.sys_id_reset_reset_bridge_in_reset_reset                              (rst_controller_reset_out_reset),                                         //                              sys_id_reset_reset_bridge_in_reset.reset
		.pixel_clk_pll_reconfig_mgmt_avalon_slave_address                      (mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_address),     //                        pixel_clk_pll_reconfig_mgmt_avalon_slave.address
		.pixel_clk_pll_reconfig_mgmt_avalon_slave_write                        (mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_write),       //                                                                .write
		.pixel_clk_pll_reconfig_mgmt_avalon_slave_read                         (mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_read),        //                                                                .read
		.pixel_clk_pll_reconfig_mgmt_avalon_slave_readdata                     (mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_readdata),    //                                                                .readdata
		.pixel_clk_pll_reconfig_mgmt_avalon_slave_writedata                    (mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_writedata),   //                                                                .writedata
		.pixel_clk_pll_reconfig_mgmt_avalon_slave_waitrequest                  (mm_interconnect_1_pixel_clk_pll_reconfig_mgmt_avalon_slave_waitrequest), //                                                                .waitrequest
		.sys_gpio_bd_s1_address                                                (mm_interconnect_1_sys_gpio_bd_s1_address),                               //                                                  sys_gpio_bd_s1.address
		.sys_gpio_bd_s1_write                                                  (mm_interconnect_1_sys_gpio_bd_s1_write),                                 //                                                                .write
		.sys_gpio_bd_s1_readdata                                               (mm_interconnect_1_sys_gpio_bd_s1_readdata),                              //                                                                .readdata
		.sys_gpio_bd_s1_writedata                                              (mm_interconnect_1_sys_gpio_bd_s1_writedata),                             //                                                                .writedata
		.sys_gpio_bd_s1_chipselect                                             (mm_interconnect_1_sys_gpio_bd_s1_chipselect),                            //                                                                .chipselect
		.sys_gpio_in_s1_address                                                (mm_interconnect_1_sys_gpio_in_s1_address),                               //                                                  sys_gpio_in_s1.address
		.sys_gpio_in_s1_write                                                  (mm_interconnect_1_sys_gpio_in_s1_write),                                 //                                                                .write
		.sys_gpio_in_s1_readdata                                               (mm_interconnect_1_sys_gpio_in_s1_readdata),                              //                                                                .readdata
		.sys_gpio_in_s1_writedata                                              (mm_interconnect_1_sys_gpio_in_s1_writedata),                             //                                                                .writedata
		.sys_gpio_in_s1_chipselect                                             (mm_interconnect_1_sys_gpio_in_s1_chipselect),                            //                                                                .chipselect
		.sys_gpio_out_s1_address                                               (mm_interconnect_1_sys_gpio_out_s1_address),                              //                                                 sys_gpio_out_s1.address
		.sys_gpio_out_s1_write                                                 (mm_interconnect_1_sys_gpio_out_s1_write),                                //                                                                .write
		.sys_gpio_out_s1_readdata                                              (mm_interconnect_1_sys_gpio_out_s1_readdata),                             //                                                                .readdata
		.sys_gpio_out_s1_writedata                                             (mm_interconnect_1_sys_gpio_out_s1_writedata),                            //                                                                .writedata
		.sys_gpio_out_s1_chipselect                                            (mm_interconnect_1_sys_gpio_out_s1_chipselect),                           //                                                                .chipselect
		.sys_id_control_slave_address                                          (mm_interconnect_1_sys_id_control_slave_address),                         //                                            sys_id_control_slave.address
		.sys_id_control_slave_readdata                                         (mm_interconnect_1_sys_id_control_slave_readdata),                        //                                                                .readdata
		.sys_spi_spi_control_port_address                                      (mm_interconnect_1_sys_spi_spi_control_port_address),                     //                                        sys_spi_spi_control_port.address
		.sys_spi_spi_control_port_write                                        (mm_interconnect_1_sys_spi_spi_control_port_write),                       //                                                                .write
		.sys_spi_spi_control_port_read                                         (mm_interconnect_1_sys_spi_spi_control_port_read),                        //                                                                .read
		.sys_spi_spi_control_port_readdata                                     (mm_interconnect_1_sys_spi_spi_control_port_readdata),                    //                                                                .readdata
		.sys_spi_spi_control_port_writedata                                    (mm_interconnect_1_sys_spi_spi_control_port_writedata),                   //                                                                .writedata
		.sys_spi_spi_control_port_chipselect                                   (mm_interconnect_1_sys_spi_spi_control_port_chipselect)                   //                                                                .chipselect
	);

	system_bd_mm_interconnect_2 mm_interconnect_2 (
		.axi_adc_dma_m_dest_axi_awid                                          (axi_adc_dma_m_dest_axi_awid),                       //                                         axi_adc_dma_m_dest_axi.awid
		.axi_adc_dma_m_dest_axi_awaddr                                        (axi_adc_dma_m_dest_axi_awaddr),                     //                                                               .awaddr
		.axi_adc_dma_m_dest_axi_awlen                                         (axi_adc_dma_m_dest_axi_awlen),                      //                                                               .awlen
		.axi_adc_dma_m_dest_axi_awsize                                        (axi_adc_dma_m_dest_axi_awsize),                     //                                                               .awsize
		.axi_adc_dma_m_dest_axi_awburst                                       (axi_adc_dma_m_dest_axi_awburst),                    //                                                               .awburst
		.axi_adc_dma_m_dest_axi_awlock                                        (axi_adc_dma_m_dest_axi_awlock),                     //                                                               .awlock
		.axi_adc_dma_m_dest_axi_awcache                                       (axi_adc_dma_m_dest_axi_awcache),                    //                                                               .awcache
		.axi_adc_dma_m_dest_axi_awprot                                        (axi_adc_dma_m_dest_axi_awprot),                     //                                                               .awprot
		.axi_adc_dma_m_dest_axi_awvalid                                       (axi_adc_dma_m_dest_axi_awvalid),                    //                                                               .awvalid
		.axi_adc_dma_m_dest_axi_awready                                       (axi_adc_dma_m_dest_axi_awready),                    //                                                               .awready
		.axi_adc_dma_m_dest_axi_wid                                           (axi_adc_dma_m_dest_axi_wid),                        //                                                               .wid
		.axi_adc_dma_m_dest_axi_wdata                                         (axi_adc_dma_m_dest_axi_wdata),                      //                                                               .wdata
		.axi_adc_dma_m_dest_axi_wstrb                                         (axi_adc_dma_m_dest_axi_wstrb),                      //                                                               .wstrb
		.axi_adc_dma_m_dest_axi_wlast                                         (axi_adc_dma_m_dest_axi_wlast),                      //                                                               .wlast
		.axi_adc_dma_m_dest_axi_wvalid                                        (axi_adc_dma_m_dest_axi_wvalid),                     //                                                               .wvalid
		.axi_adc_dma_m_dest_axi_wready                                        (axi_adc_dma_m_dest_axi_wready),                     //                                                               .wready
		.axi_adc_dma_m_dest_axi_bid                                           (axi_adc_dma_m_dest_axi_bid),                        //                                                               .bid
		.axi_adc_dma_m_dest_axi_bresp                                         (axi_adc_dma_m_dest_axi_bresp),                      //                                                               .bresp
		.axi_adc_dma_m_dest_axi_bvalid                                        (axi_adc_dma_m_dest_axi_bvalid),                     //                                                               .bvalid
		.axi_adc_dma_m_dest_axi_bready                                        (axi_adc_dma_m_dest_axi_bready),                     //                                                               .bready
		.axi_adc_dma_m_dest_axi_arid                                          (axi_adc_dma_m_dest_axi_arid),                       //                                                               .arid
		.axi_adc_dma_m_dest_axi_araddr                                        (axi_adc_dma_m_dest_axi_araddr),                     //                                                               .araddr
		.axi_adc_dma_m_dest_axi_arlen                                         (axi_adc_dma_m_dest_axi_arlen),                      //                                                               .arlen
		.axi_adc_dma_m_dest_axi_arsize                                        (axi_adc_dma_m_dest_axi_arsize),                     //                                                               .arsize
		.axi_adc_dma_m_dest_axi_arburst                                       (axi_adc_dma_m_dest_axi_arburst),                    //                                                               .arburst
		.axi_adc_dma_m_dest_axi_arlock                                        (axi_adc_dma_m_dest_axi_arlock),                     //                                                               .arlock
		.axi_adc_dma_m_dest_axi_arcache                                       (axi_adc_dma_m_dest_axi_arcache),                    //                                                               .arcache
		.axi_adc_dma_m_dest_axi_arprot                                        (axi_adc_dma_m_dest_axi_arprot),                     //                                                               .arprot
		.axi_adc_dma_m_dest_axi_arvalid                                       (axi_adc_dma_m_dest_axi_arvalid),                    //                                                               .arvalid
		.axi_adc_dma_m_dest_axi_arready                                       (axi_adc_dma_m_dest_axi_arready),                    //                                                               .arready
		.axi_adc_dma_m_dest_axi_rid                                           (axi_adc_dma_m_dest_axi_rid),                        //                                                               .rid
		.axi_adc_dma_m_dest_axi_rdata                                         (axi_adc_dma_m_dest_axi_rdata),                      //                                                               .rdata
		.axi_adc_dma_m_dest_axi_rresp                                         (axi_adc_dma_m_dest_axi_rresp),                      //                                                               .rresp
		.axi_adc_dma_m_dest_axi_rlast                                         (axi_adc_dma_m_dest_axi_rlast),                      //                                                               .rlast
		.axi_adc_dma_m_dest_axi_rvalid                                        (axi_adc_dma_m_dest_axi_rvalid),                     //                                                               .rvalid
		.axi_adc_dma_m_dest_axi_rready                                        (axi_adc_dma_m_dest_axi_rready),                     //                                                               .rready
		.sys_hps_f2h_sdram1_data_awid                                         (mm_interconnect_2_sys_hps_f2h_sdram1_data_awid),    //                                        sys_hps_f2h_sdram1_data.awid
		.sys_hps_f2h_sdram1_data_awaddr                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_awaddr),  //                                                               .awaddr
		.sys_hps_f2h_sdram1_data_awlen                                        (mm_interconnect_2_sys_hps_f2h_sdram1_data_awlen),   //                                                               .awlen
		.sys_hps_f2h_sdram1_data_awsize                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_awsize),  //                                                               .awsize
		.sys_hps_f2h_sdram1_data_awburst                                      (mm_interconnect_2_sys_hps_f2h_sdram1_data_awburst), //                                                               .awburst
		.sys_hps_f2h_sdram1_data_awlock                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_awlock),  //                                                               .awlock
		.sys_hps_f2h_sdram1_data_awcache                                      (mm_interconnect_2_sys_hps_f2h_sdram1_data_awcache), //                                                               .awcache
		.sys_hps_f2h_sdram1_data_awprot                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_awprot),  //                                                               .awprot
		.sys_hps_f2h_sdram1_data_awvalid                                      (mm_interconnect_2_sys_hps_f2h_sdram1_data_awvalid), //                                                               .awvalid
		.sys_hps_f2h_sdram1_data_awready                                      (mm_interconnect_2_sys_hps_f2h_sdram1_data_awready), //                                                               .awready
		.sys_hps_f2h_sdram1_data_wid                                          (mm_interconnect_2_sys_hps_f2h_sdram1_data_wid),     //                                                               .wid
		.sys_hps_f2h_sdram1_data_wdata                                        (mm_interconnect_2_sys_hps_f2h_sdram1_data_wdata),   //                                                               .wdata
		.sys_hps_f2h_sdram1_data_wstrb                                        (mm_interconnect_2_sys_hps_f2h_sdram1_data_wstrb),   //                                                               .wstrb
		.sys_hps_f2h_sdram1_data_wlast                                        (mm_interconnect_2_sys_hps_f2h_sdram1_data_wlast),   //                                                               .wlast
		.sys_hps_f2h_sdram1_data_wvalid                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_wvalid),  //                                                               .wvalid
		.sys_hps_f2h_sdram1_data_wready                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_wready),  //                                                               .wready
		.sys_hps_f2h_sdram1_data_bid                                          (mm_interconnect_2_sys_hps_f2h_sdram1_data_bid),     //                                                               .bid
		.sys_hps_f2h_sdram1_data_bresp                                        (mm_interconnect_2_sys_hps_f2h_sdram1_data_bresp),   //                                                               .bresp
		.sys_hps_f2h_sdram1_data_bvalid                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_bvalid),  //                                                               .bvalid
		.sys_hps_f2h_sdram1_data_bready                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_bready),  //                                                               .bready
		.sys_hps_f2h_sdram1_data_arid                                         (mm_interconnect_2_sys_hps_f2h_sdram1_data_arid),    //                                                               .arid
		.sys_hps_f2h_sdram1_data_araddr                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_araddr),  //                                                               .araddr
		.sys_hps_f2h_sdram1_data_arlen                                        (mm_interconnect_2_sys_hps_f2h_sdram1_data_arlen),   //                                                               .arlen
		.sys_hps_f2h_sdram1_data_arsize                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_arsize),  //                                                               .arsize
		.sys_hps_f2h_sdram1_data_arburst                                      (mm_interconnect_2_sys_hps_f2h_sdram1_data_arburst), //                                                               .arburst
		.sys_hps_f2h_sdram1_data_arlock                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_arlock),  //                                                               .arlock
		.sys_hps_f2h_sdram1_data_arcache                                      (mm_interconnect_2_sys_hps_f2h_sdram1_data_arcache), //                                                               .arcache
		.sys_hps_f2h_sdram1_data_arprot                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_arprot),  //                                                               .arprot
		.sys_hps_f2h_sdram1_data_arvalid                                      (mm_interconnect_2_sys_hps_f2h_sdram1_data_arvalid), //                                                               .arvalid
		.sys_hps_f2h_sdram1_data_arready                                      (mm_interconnect_2_sys_hps_f2h_sdram1_data_arready), //                                                               .arready
		.sys_hps_f2h_sdram1_data_rid                                          (mm_interconnect_2_sys_hps_f2h_sdram1_data_rid),     //                                                               .rid
		.sys_hps_f2h_sdram1_data_rdata                                        (mm_interconnect_2_sys_hps_f2h_sdram1_data_rdata),   //                                                               .rdata
		.sys_hps_f2h_sdram1_data_rresp                                        (mm_interconnect_2_sys_hps_f2h_sdram1_data_rresp),   //                                                               .rresp
		.sys_hps_f2h_sdram1_data_rlast                                        (mm_interconnect_2_sys_hps_f2h_sdram1_data_rlast),   //                                                               .rlast
		.sys_hps_f2h_sdram1_data_rvalid                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_rvalid),  //                                                               .rvalid
		.sys_hps_f2h_sdram1_data_rready                                       (mm_interconnect_2_sys_hps_f2h_sdram1_data_rready),  //                                                               .rready
		.sys_clk_clk_clk                                                      (sys_clk_clk),                                       //                                                    sys_clk_clk.clk
		.sys_dma_clk_clk_clk                                                  (sys_hps_h2f_user0_clock_clk),                       //                                                sys_dma_clk_clk.clk
		.axi_adc_dma_m_dest_axi_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                    //             axi_adc_dma_m_dest_axi_reset_reset_bridge_in_reset.reset
		.sys_hps_f2h_sdram1_data_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset)                 // sys_hps_f2h_sdram1_data_agent_reset_sink_reset_bridge_in_reset.reset
	);

	system_bd_mm_interconnect_3 mm_interconnect_3 (
		.sys_hps_f2h_sdram0_data_awid                                      (mm_interconnect_3_sys_hps_f2h_sdram0_data_awid),    //                                     sys_hps_f2h_sdram0_data.awid
		.sys_hps_f2h_sdram0_data_awaddr                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_awaddr),  //                                                            .awaddr
		.sys_hps_f2h_sdram0_data_awlen                                     (mm_interconnect_3_sys_hps_f2h_sdram0_data_awlen),   //                                                            .awlen
		.sys_hps_f2h_sdram0_data_awsize                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_awsize),  //                                                            .awsize
		.sys_hps_f2h_sdram0_data_awburst                                   (mm_interconnect_3_sys_hps_f2h_sdram0_data_awburst), //                                                            .awburst
		.sys_hps_f2h_sdram0_data_awlock                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_awlock),  //                                                            .awlock
		.sys_hps_f2h_sdram0_data_awcache                                   (mm_interconnect_3_sys_hps_f2h_sdram0_data_awcache), //                                                            .awcache
		.sys_hps_f2h_sdram0_data_awprot                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_awprot),  //                                                            .awprot
		.sys_hps_f2h_sdram0_data_awvalid                                   (mm_interconnect_3_sys_hps_f2h_sdram0_data_awvalid), //                                                            .awvalid
		.sys_hps_f2h_sdram0_data_awready                                   (mm_interconnect_3_sys_hps_f2h_sdram0_data_awready), //                                                            .awready
		.sys_hps_f2h_sdram0_data_wid                                       (mm_interconnect_3_sys_hps_f2h_sdram0_data_wid),     //                                                            .wid
		.sys_hps_f2h_sdram0_data_wdata                                     (mm_interconnect_3_sys_hps_f2h_sdram0_data_wdata),   //                                                            .wdata
		.sys_hps_f2h_sdram0_data_wstrb                                     (mm_interconnect_3_sys_hps_f2h_sdram0_data_wstrb),   //                                                            .wstrb
		.sys_hps_f2h_sdram0_data_wlast                                     (mm_interconnect_3_sys_hps_f2h_sdram0_data_wlast),   //                                                            .wlast
		.sys_hps_f2h_sdram0_data_wvalid                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_wvalid),  //                                                            .wvalid
		.sys_hps_f2h_sdram0_data_wready                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_wready),  //                                                            .wready
		.sys_hps_f2h_sdram0_data_bid                                       (mm_interconnect_3_sys_hps_f2h_sdram0_data_bid),     //                                                            .bid
		.sys_hps_f2h_sdram0_data_bresp                                     (mm_interconnect_3_sys_hps_f2h_sdram0_data_bresp),   //                                                            .bresp
		.sys_hps_f2h_sdram0_data_bvalid                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_bvalid),  //                                                            .bvalid
		.sys_hps_f2h_sdram0_data_bready                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_bready),  //                                                            .bready
		.sys_hps_f2h_sdram0_data_arid                                      (mm_interconnect_3_sys_hps_f2h_sdram0_data_arid),    //                                                            .arid
		.sys_hps_f2h_sdram0_data_araddr                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_araddr),  //                                                            .araddr
		.sys_hps_f2h_sdram0_data_arlen                                     (mm_interconnect_3_sys_hps_f2h_sdram0_data_arlen),   //                                                            .arlen
		.sys_hps_f2h_sdram0_data_arsize                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_arsize),  //                                                            .arsize
		.sys_hps_f2h_sdram0_data_arburst                                   (mm_interconnect_3_sys_hps_f2h_sdram0_data_arburst), //                                                            .arburst
		.sys_hps_f2h_sdram0_data_arlock                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_arlock),  //                                                            .arlock
		.sys_hps_f2h_sdram0_data_arcache                                   (mm_interconnect_3_sys_hps_f2h_sdram0_data_arcache), //                                                            .arcache
		.sys_hps_f2h_sdram0_data_arprot                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_arprot),  //                                                            .arprot
		.sys_hps_f2h_sdram0_data_arvalid                                   (mm_interconnect_3_sys_hps_f2h_sdram0_data_arvalid), //                                                            .arvalid
		.sys_hps_f2h_sdram0_data_arready                                   (mm_interconnect_3_sys_hps_f2h_sdram0_data_arready), //                                                            .arready
		.sys_hps_f2h_sdram0_data_rid                                       (mm_interconnect_3_sys_hps_f2h_sdram0_data_rid),     //                                                            .rid
		.sys_hps_f2h_sdram0_data_rdata                                     (mm_interconnect_3_sys_hps_f2h_sdram0_data_rdata),   //                                                            .rdata
		.sys_hps_f2h_sdram0_data_rresp                                     (mm_interconnect_3_sys_hps_f2h_sdram0_data_rresp),   //                                                            .rresp
		.sys_hps_f2h_sdram0_data_rlast                                     (mm_interconnect_3_sys_hps_f2h_sdram0_data_rlast),   //                                                            .rlast
		.sys_hps_f2h_sdram0_data_rvalid                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_rvalid),  //                                                            .rvalid
		.sys_hps_f2h_sdram0_data_rready                                    (mm_interconnect_3_sys_hps_f2h_sdram0_data_rready),  //                                                            .rready
		.video_dmac_m_src_axi_awid                                         (video_dmac_m_src_axi_awid),                         //                                        video_dmac_m_src_axi.awid
		.video_dmac_m_src_axi_awaddr                                       (video_dmac_m_src_axi_awaddr),                       //                                                            .awaddr
		.video_dmac_m_src_axi_awlen                                        (video_dmac_m_src_axi_awlen),                        //                                                            .awlen
		.video_dmac_m_src_axi_awsize                                       (video_dmac_m_src_axi_awsize),                       //                                                            .awsize
		.video_dmac_m_src_axi_awburst                                      (video_dmac_m_src_axi_awburst),                      //                                                            .awburst
		.video_dmac_m_src_axi_awlock                                       (video_dmac_m_src_axi_awlock),                       //                                                            .awlock
		.video_dmac_m_src_axi_awcache                                      (video_dmac_m_src_axi_awcache),                      //                                                            .awcache
		.video_dmac_m_src_axi_awprot                                       (video_dmac_m_src_axi_awprot),                       //                                                            .awprot
		.video_dmac_m_src_axi_awvalid                                      (video_dmac_m_src_axi_awvalid),                      //                                                            .awvalid
		.video_dmac_m_src_axi_awready                                      (video_dmac_m_src_axi_awready),                      //                                                            .awready
		.video_dmac_m_src_axi_wid                                          (video_dmac_m_src_axi_wid),                          //                                                            .wid
		.video_dmac_m_src_axi_wdata                                        (video_dmac_m_src_axi_wdata),                        //                                                            .wdata
		.video_dmac_m_src_axi_wstrb                                        (video_dmac_m_src_axi_wstrb),                        //                                                            .wstrb
		.video_dmac_m_src_axi_wlast                                        (video_dmac_m_src_axi_wlast),                        //                                                            .wlast
		.video_dmac_m_src_axi_wvalid                                       (video_dmac_m_src_axi_wvalid),                       //                                                            .wvalid
		.video_dmac_m_src_axi_wready                                       (video_dmac_m_src_axi_wready),                       //                                                            .wready
		.video_dmac_m_src_axi_bid                                          (video_dmac_m_src_axi_bid),                          //                                                            .bid
		.video_dmac_m_src_axi_bresp                                        (video_dmac_m_src_axi_bresp),                        //                                                            .bresp
		.video_dmac_m_src_axi_bvalid                                       (video_dmac_m_src_axi_bvalid),                       //                                                            .bvalid
		.video_dmac_m_src_axi_bready                                       (video_dmac_m_src_axi_bready),                       //                                                            .bready
		.video_dmac_m_src_axi_arid                                         (video_dmac_m_src_axi_arid),                         //                                                            .arid
		.video_dmac_m_src_axi_araddr                                       (video_dmac_m_src_axi_araddr),                       //                                                            .araddr
		.video_dmac_m_src_axi_arlen                                        (video_dmac_m_src_axi_arlen),                        //                                                            .arlen
		.video_dmac_m_src_axi_arsize                                       (video_dmac_m_src_axi_arsize),                       //                                                            .arsize
		.video_dmac_m_src_axi_arburst                                      (video_dmac_m_src_axi_arburst),                      //                                                            .arburst
		.video_dmac_m_src_axi_arlock                                       (video_dmac_m_src_axi_arlock),                       //                                                            .arlock
		.video_dmac_m_src_axi_arcache                                      (video_dmac_m_src_axi_arcache),                      //                                                            .arcache
		.video_dmac_m_src_axi_arprot                                       (video_dmac_m_src_axi_arprot),                       //                                                            .arprot
		.video_dmac_m_src_axi_arvalid                                      (video_dmac_m_src_axi_arvalid),                      //                                                            .arvalid
		.video_dmac_m_src_axi_arready                                      (video_dmac_m_src_axi_arready),                      //                                                            .arready
		.video_dmac_m_src_axi_rid                                          (video_dmac_m_src_axi_rid),                          //                                                            .rid
		.video_dmac_m_src_axi_rdata                                        (video_dmac_m_src_axi_rdata),                        //                                                            .rdata
		.video_dmac_m_src_axi_rresp                                        (video_dmac_m_src_axi_rresp),                        //                                                            .rresp
		.video_dmac_m_src_axi_rlast                                        (video_dmac_m_src_axi_rlast),                        //                                                            .rlast
		.video_dmac_m_src_axi_rvalid                                       (video_dmac_m_src_axi_rvalid),                       //                                                            .rvalid
		.video_dmac_m_src_axi_rready                                       (video_dmac_m_src_axi_rready),                       //                                                            .rready
		.pixel_clk_pll_outclk1_clk                                         (pixel_clk_pll_outclk1_clk),                         //                                       pixel_clk_pll_outclk1.clk
		.video_dmac_m_src_axi_id_pad_clk_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                // video_dmac_m_src_axi_id_pad_clk_reset_reset_bridge_in_reset.reset
		.video_dmac_m_src_axi_reset_reset_bridge_in_reset_reset            (rst_controller_001_reset_out_reset)                 //            video_dmac_m_src_axi_reset_reset_bridge_in_reset.reset
	);

	system_bd_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq), // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq), // receiver3.irq
		.sender_irq    (sys_hps_f2h_irq0_irq)      //    sender.irq
	);

	system_bd_irq_mapper_001 irq_mapper_001 (
		.clk        (),                     //       clk.clk
		.reset      (),                     // clk_reset.reset
		.sender_irq (sys_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~sys_rst_reset_n),                   // reset_in0.reset
		.clk            (sys_clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~sys_rst_reset_n),                   // reset_in0.reset
		.clk            (pixel_clk_pll_outclk1_clk),          //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~sys_hps_h2f_reset_reset_n),         // reset_in0.reset
		.clk            (sys_clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~sys_hps_h2f_reset_reset_n),         // reset_in0.reset
		.clk            (sys_hps_h2f_user0_clock_clk),        //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~sys_hps_h2f_reset_reset_n),         // reset_in0.reset
		.clk            (pixel_clk_pll_outclk1_clk),          //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
